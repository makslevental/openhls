module fsqrt#(parameter ID=1)
  (input  clk,
   input  [16:0] X,
   output [16:0] R);
  wire [6:0] fracx;
  wire [6:0] ern0;
  wire [2:0] xsx;
  wire [6:0] ern1;
  wire [6:0] ern1_d1;
  wire [6:0] ern1_d2;
  wire [10:0] fracxnorm;
  wire [1:0] s0;
  wire [10:0] t1;
  wire d1;
  wire [11:0] t1s;
  wire [5:0] t1s_h;
  wire [5:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [10:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [11:0] t2s;
  wire [6:0] t2s_h;
  wire [4:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [10:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [11:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [3:0] t3s_l;
  wire [3:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [10:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [11:0] t4s;
  wire [8:0] t4s_h;
  wire [2:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [10:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [11:0] t5s;
  wire [9:0] t5s_h;
  wire [1:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [10:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [11:0] t6s;
  wire [10:0] t6s_h;
  wire t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [10:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [11:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [10:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d9;
  wire [9:0] mr;
  wire [6:0] fr;
  wire round;
  wire [6:0] frrnd;
  wire [13:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [6:0] n18_o;
  wire [5:0] n19_o;
  wire [6:0] n21_o;
  wire [2:0] n22_o;
  wire [6:0] n24_o;
  wire n25_o;
  wire [6:0] n26_o;
  wire [6:0] n27_o;
  wire [7:0] n29_o;
  wire [10:0] n31_o;
  wire n32_o;
  wire n33_o;
  wire [10:0] n34_o;
  wire [8:0] n36_o;
  wire [10:0] n38_o;
  wire [3:0] n40_o;
  wire [3:0] n42_o;
  wire [6:0] n43_o;
  wire [10:0] n44_o;
  wire n45_o;
  wire n46_o;
  wire [11:0] n48_o;
  wire [5:0] n49_o;
  wire [5:0] n50_o;
  wire [2:0] n52_o;
  wire [3:0] n53_o;
  wire n54_o;
  wire [4:0] n55_o;
  wire [5:0] n57_o;
  wire [5:0] n58_o;
  wire [5:0] n59_o;
  wire [5:0] n60_o;
  wire [4:0] n61_o;
  wire [10:0] n62_o;
  wire [2:0] n63_o;
  wire n64_o;
  wire n65_o;
  wire [11:0] n67_o;
  wire [6:0] n68_o;
  wire [4:0] n69_o;
  wire [3:0] n71_o;
  wire [4:0] n72_o;
  wire n73_o;
  wire [5:0] n74_o;
  wire [6:0] n76_o;
  wire [6:0] n77_o;
  wire [6:0] n78_o;
  wire [6:0] n79_o;
  wire [5:0] n80_o;
  wire [10:0] n81_o;
  wire [3:0] n82_o;
  wire n83_o;
  wire n84_o;
  wire [11:0] n86_o;
  wire [7:0] n87_o;
  wire [3:0] n88_o;
  wire [4:0] n90_o;
  wire [5:0] n91_o;
  wire n92_o;
  wire [6:0] n93_o;
  wire [7:0] n95_o;
  wire [7:0] n96_o;
  wire [7:0] n97_o;
  wire [7:0] n98_o;
  wire [6:0] n99_o;
  wire [10:0] n100_o;
  wire [4:0] n101_o;
  wire n102_o;
  wire n103_o;
  wire [11:0] n105_o;
  wire [8:0] n106_o;
  wire [2:0] n107_o;
  wire [5:0] n109_o;
  wire [6:0] n110_o;
  wire n111_o;
  wire [7:0] n112_o;
  wire [8:0] n114_o;
  wire [8:0] n115_o;
  wire [8:0] n116_o;
  wire [8:0] n117_o;
  wire [7:0] n118_o;
  wire [10:0] n119_o;
  wire [5:0] n120_o;
  wire n121_o;
  wire n122_o;
  wire [11:0] n124_o;
  wire [9:0] n125_o;
  wire [1:0] n126_o;
  wire [6:0] n128_o;
  wire [7:0] n129_o;
  wire n130_o;
  wire [8:0] n131_o;
  wire [9:0] n133_o;
  wire [9:0] n134_o;
  wire [9:0] n135_o;
  wire [9:0] n136_o;
  wire [8:0] n137_o;
  wire [10:0] n138_o;
  wire [6:0] n139_o;
  wire n140_o;
  wire n141_o;
  wire [11:0] n143_o;
  wire [10:0] n144_o;
  wire n145_o;
  wire [7:0] n147_o;
  wire [8:0] n148_o;
  wire n149_o;
  wire [9:0] n150_o;
  wire [10:0] n152_o;
  wire [10:0] n153_o;
  wire [10:0] n154_o;
  wire [10:0] n155_o;
  wire [9:0] n156_o;
  wire [10:0] n157_o;
  wire [7:0] n158_o;
  wire n159_o;
  wire n160_o;
  wire [11:0] n162_o;
  wire [8:0] n164_o;
  wire [9:0] n165_o;
  wire n166_o;
  wire [10:0] n167_o;
  wire [11:0] n169_o;
  wire [11:0] n170_o;
  wire [11:0] n171_o;
  wire [11:0] n172_o;
  wire [10:0] n173_o;
  wire [8:0] n174_o;
  wire n175_o;
  wire n176_o;
  wire [9:0] n177_o;
  wire [6:0] n178_o;
  wire n179_o;
  wire [6:0] n181_o;
  wire [6:0] n182_o;
  wire [13:0] n183_o;
  wire n186_o;
  wire n189_o;
  wire n192_o;
  wire n195_o;
  wire [3:0] n197_o;
  reg [2:0] n198_o;
  wire [16:0] n199_o;
  reg [6:0] n200_q;
  reg [6:0] n201_q;
  reg n202_q;
  reg [7:0] n203_q;
  reg [3:0] n204_q;
  reg [7:0] n205_q;
  reg [4:0] n206_q;
  reg n207_q;
  reg [11:0] n208_q;
  reg [11:0] n209_q;
  reg [8:0] n210_q;
  reg [2:0] n211_q;
  reg [2:0] n212_q;
  assign R = n199_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:30:8  */
  assign fracx = n18_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:31:8  */
  assign ern0 = n21_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:32:8  */
  assign xsx = n22_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:33:8  */
  assign ern1 = n27_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:33:14  */
  assign ern1_d1 = n200_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:33:23  */
  assign ern1_d2 = n201_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:34:8  */
  assign fracxnorm = n34_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:36:8  */
  assign t1 = n44_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:37:8  */
  assign d1 = n46_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:38:8  */
  assign t1s = n48_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:39:8  */
  assign t1s_h = n49_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:40:8  */
  assign t1s_l = n50_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:41:8  */
  assign u1 = n57_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:42:8  */
  assign t3_h = n59_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:43:8  */
  assign t2 = n62_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:44:8  */
  assign s1 = n63_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:45:8  */
  assign d2 = n65_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:46:8  */
  assign t2s = n67_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:47:8  */
  assign t2s_h = n68_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:48:8  */
  assign t2s_l = n69_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:49:8  */
  assign u2 = n76_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:50:8  */
  assign t4_h = n78_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:51:8  */
  assign t3 = n81_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:52:8  */
  assign s2 = n82_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:53:8  */
  assign d3 = n84_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:53:12  */
  assign d3_d1 = n202_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:54:8  */
  assign t3s = n86_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:55:8  */
  assign t3s_h = n87_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:55:15  */
  assign t3s_h_d1 = n203_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:56:8  */
  assign t3s_l = n88_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:56:15  */
  assign t3s_l_d1 = n204_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:57:8  */
  assign u3 = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:57:12  */
  assign u3_d1 = n205_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:58:8  */
  assign t5_h = n97_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:59:8  */
  assign t4 = n100_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:60:8  */
  assign s3 = n101_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:60:12  */
  assign s3_d1 = n206_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:61:8  */
  assign d4 = n103_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:62:8  */
  assign t4s = n105_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:63:8  */
  assign t4s_h = n106_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:64:8  */
  assign t4s_l = n107_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:65:8  */
  assign u4 = n114_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:66:8  */
  assign t6_h = n116_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:67:8  */
  assign t5 = n119_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:68:8  */
  assign s4 = n120_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:69:8  */
  assign d5 = n122_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:70:8  */
  assign t5s = n124_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:71:8  */
  assign t5s_h = n125_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:72:8  */
  assign t5s_l = n126_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:73:8  */
  assign u5 = n133_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:74:8  */
  assign t7_h = n135_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:75:8  */
  assign t6 = n138_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:76:8  */
  assign s5 = n139_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:77:8  */
  assign d6 = n141_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:78:8  */
  assign t6s = n143_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:79:8  */
  assign t6s_h = n144_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:80:8  */
  assign t6s_l = n145_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:81:8  */
  assign u6 = n152_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:82:8  */
  assign t8_h = n154_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:83:8  */
  assign t7 = n157_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:84:8  */
  assign s6 = n158_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:85:8  */
  assign d7 = n160_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:85:12  */
  assign d7_d1 = n207_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:191:16  */
  assign t7s = n162_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:87:8  */
  assign t7s_h = t7s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:87:15  */
  assign t7s_h_d1 = n208_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:88:8  */
  assign u7 = n169_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:88:12  */
  assign u7_d1 = n209_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:89:8  */
  assign t9_h = n171_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:90:8  */
  assign t8 = n173_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:91:8  */
  assign s7 = n174_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:91:12  */
  assign s7_d1 = n210_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:92:8  */
  assign d9 = n176_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:93:8  */
  assign mr = n177_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:94:8  */
  assign fr = n178_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:95:8  */
  assign round = n179_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:96:8  */
  assign frrnd = n182_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:97:8  */
  assign rn2 = n183_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:98:8  */
  assign xsr = n198_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:98:13  */
  assign xsr_d1 = n211_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:98:21  */
  assign xsr_d2 = n212_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:118:14  */
  assign n18_o = X[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:119:19  */
  assign n19_o = X[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:119:16  */
  assign n21_o = {1'b0, n19_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:120:12  */
  assign n22_o = X[16:14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:121:17  */
  assign n24_o = ern0 + 7'b0011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:121:51  */
  assign n25_o = X[7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:121:48  */
  assign n26_o = {6'b0, n25_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:121:48  */
  assign n27_o = n24_o + n26_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:122:21  */
  assign n29_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:122:29  */
  assign n31_o = {n29_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:122:43  */
  assign n32_o = X[7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:122:47  */
  assign n33_o = ~n32_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:122:37  */
  assign n34_o = n33_o ? n31_o : n38_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:123:15  */
  assign n36_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:123:22  */
  assign n38_o = {n36_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:125:29  */
  assign n40_o = fracxnorm[10:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:125:18  */
  assign n42_o = 4'b0111 + n40_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:125:55  */
  assign n43_o = fracxnorm[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:125:44  */
  assign n44_o = {n42_o, n43_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:129:16  */
  assign n45_o = t1[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:129:10  */
  assign n46_o = ~n45_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:130:14  */
  assign n48_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:131:16  */
  assign n49_o = t1s[11:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:132:16  */
  assign n50_o = t1s[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:133:15  */
  assign n52_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:133:20  */
  assign n53_o = {n52_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:133:28  */
  assign n54_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:133:25  */
  assign n55_o = {n53_o, n54_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:133:36  */
  assign n57_o = {n55_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:134:20  */
  assign n58_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:134:25  */
  assign n59_o = d1 ? n58_o : n60_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:135:20  */
  assign n60_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:136:14  */
  assign n61_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:136:27  */
  assign n62_o = {n61_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:137:13  */
  assign n63_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:139:16  */
  assign n64_o = t2[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:139:10  */
  assign n65_o = ~n64_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:140:14  */
  assign n67_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:141:16  */
  assign n68_o = t2s[11:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:142:16  */
  assign n69_o = t2s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:143:15  */
  assign n71_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:143:20  */
  assign n72_o = {n71_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:143:28  */
  assign n73_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:143:25  */
  assign n74_o = {n72_o, n73_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:143:36  */
  assign n76_o = {n74_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:144:20  */
  assign n77_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:144:25  */
  assign n78_o = d2 ? n77_o : n79_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:145:20  */
  assign n79_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:146:14  */
  assign n80_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:146:27  */
  assign n81_o = {n80_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:147:13  */
  assign n82_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:149:16  */
  assign n83_o = t3[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:149:10  */
  assign n84_o = ~n83_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:150:14  */
  assign n86_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:151:16  */
  assign n87_o = t3s[11:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:152:16  */
  assign n88_o = t3s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:153:15  */
  assign n90_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:153:20  */
  assign n91_o = {n90_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:153:28  */
  assign n92_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:153:25  */
  assign n93_o = {n91_o, n92_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:153:36  */
  assign n95_o = {n93_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:154:23  */
  assign n96_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:154:31  */
  assign n97_o = d3_d1 ? n96_o : n98_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:155:23  */
  assign n98_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:156:14  */
  assign n99_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:156:27  */
  assign n100_o = {n99_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:157:13  */
  assign n101_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:159:16  */
  assign n102_o = t4[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:159:10  */
  assign n103_o = ~n102_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:160:14  */
  assign n105_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:161:16  */
  assign n106_o = t4s[11:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:162:16  */
  assign n107_o = t4s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:163:15  */
  assign n109_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:163:23  */
  assign n110_o = {n109_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:163:31  */
  assign n111_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:163:28  */
  assign n112_o = {n110_o, n111_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:163:39  */
  assign n114_o = {n112_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:164:20  */
  assign n115_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:164:25  */
  assign n116_o = d4 ? n115_o : n117_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:165:20  */
  assign n117_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:166:14  */
  assign n118_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:166:27  */
  assign n119_o = {n118_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:167:16  */
  assign n120_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:169:16  */
  assign n121_o = t5[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:169:10  */
  assign n122_o = ~n121_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:170:14  */
  assign n124_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:171:16  */
  assign n125_o = t5s[11:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:172:16  */
  assign n126_o = t5s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:173:15  */
  assign n128_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:173:20  */
  assign n129_o = {n128_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:173:28  */
  assign n130_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:173:25  */
  assign n131_o = {n129_o, n130_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:173:36  */
  assign n133_o = {n131_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:174:20  */
  assign n134_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:174:25  */
  assign n135_o = d5 ? n134_o : n136_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:175:20  */
  assign n136_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:176:14  */
  assign n137_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:176:27  */
  assign n138_o = {n137_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:177:13  */
  assign n139_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:179:16  */
  assign n140_o = t6[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:179:10  */
  assign n141_o = ~n140_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:180:14  */
  assign n143_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:181:16  */
  assign n144_o = t6s[11:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:182:16  */
  assign n145_o = t6s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:183:15  */
  assign n147_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:183:20  */
  assign n148_o = {n147_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:183:28  */
  assign n149_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:183:25  */
  assign n150_o = {n148_o, n149_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:183:36  */
  assign n152_o = {n150_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:184:20  */
  assign n153_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:184:25  */
  assign n154_o = d6 ? n153_o : n155_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:185:20  */
  assign n155_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:186:14  */
  assign n156_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:186:27  */
  assign n157_o = {n156_o, t6s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:187:13  */
  assign n158_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:189:16  */
  assign n159_o = t7[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:189:10  */
  assign n160_o = ~n159_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:190:14  */
  assign n162_o = {t7, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:192:15  */
  assign n164_o = {1'b0, s6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:192:20  */
  assign n165_o = {n164_o, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:192:28  */
  assign n166_o = ~d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:192:25  */
  assign n167_o = {n165_o, n166_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:192:36  */
  assign n169_o = {n167_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:193:23  */
  assign n170_o = t7s_h_d1 - u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:193:31  */
  assign n171_o = d7_d1 ? n170_o : n172_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:194:23  */
  assign n172_o = t7s_h_d1 + u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:195:14  */
  assign n173_o = t9_h[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:196:13  */
  assign n174_o = {s6, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:197:16  */
  assign n175_o = t8[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:197:10  */
  assign n176_o = ~n175_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:198:16  */
  assign n177_o = {s7_d1, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:199:12  */
  assign n178_o = mr[7:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:200:15  */
  assign n179_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:201:39  */
  assign n181_o = {6'b000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:201:16  */
  assign n182_o = fr + n181_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:202:19  */
  assign n183_o = {ern1_d2, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:205:21  */
  assign n186_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:206:21  */
  assign n189_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:207:21  */
  assign n192_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:208:21  */
  assign n195_o = xsx == 3'b001;
  assign n197_o = {n195_o, n192_o, n189_o, n186_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:204:4  */
  always @*
    case (n197_o)
      4'b1000: n198_o = 3'b001;
      4'b0100: n198_o = 3'b000;
      4'b0010: n198_o = 3'b100;
      4'b0001: n198_o = 3'b010;
      default: n198_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:210:16  */
  assign n199_o = {xsr_d2, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n200_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n201_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n202_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n203_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n204_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n205_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n206_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n207_q <= d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n208_q <= t7s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n209_q <= u7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n210_q <= s7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n211_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_7_7.vhdl:102:10  */
  always @(posedge clk)
    n212_q <= xsr_d1;
endmodule

