module fsqrt#(parameter ID=1)
  (input  clk,
   input  [18:0] X,
   output [18:0] R);
  wire [7:0] fracx;
  wire [7:0] ern0;
  wire [2:0] xsx;
  wire [7:0] ern1;
  wire [7:0] ern1_d1;
  wire [7:0] ern1_d2;
  wire [11:0] fracxnorm;
  wire [1:0] s0;
  wire [11:0] t1;
  wire d1;
  wire [12:0] t1s;
  wire [5:0] t1s_h;
  wire [6:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [11:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [12:0] t2s;
  wire [6:0] t2s_h;
  wire [5:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [11:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [12:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [4:0] t3s_l;
  wire [4:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [11:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [12:0] t4s;
  wire [8:0] t4s_h;
  wire [3:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [11:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [12:0] t5s;
  wire [9:0] t5s_h;
  wire [2:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [11:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [12:0] t6s;
  wire [10:0] t6s_h;
  wire [1:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [11:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [12:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire t7s_l;
  wire t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [11:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [12:0] t8s;
  wire [12:0] t8s_h;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [11:0] t9;
  wire [9:0] s8;
  wire d10;
  wire [10:0] mr;
  wire [7:0] fr;
  wire round;
  wire [7:0] frrnd;
  wire [15:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [7:0] n19_o;
  wire [6:0] n20_o;
  wire [7:0] n22_o;
  wire [2:0] n23_o;
  wire [7:0] n25_o;
  wire n26_o;
  wire [7:0] n27_o;
  wire [7:0] n28_o;
  wire [8:0] n30_o;
  wire [11:0] n32_o;
  wire n33_o;
  wire n34_o;
  wire [11:0] n35_o;
  wire [9:0] n37_o;
  wire [11:0] n39_o;
  wire [3:0] n41_o;
  wire [3:0] n43_o;
  wire [7:0] n44_o;
  wire [11:0] n45_o;
  wire n46_o;
  wire n47_o;
  wire [12:0] n49_o;
  wire [5:0] n50_o;
  wire [6:0] n51_o;
  wire [2:0] n53_o;
  wire [3:0] n54_o;
  wire n55_o;
  wire [4:0] n56_o;
  wire [5:0] n58_o;
  wire [5:0] n59_o;
  wire [5:0] n60_o;
  wire [5:0] n61_o;
  wire [4:0] n62_o;
  wire [11:0] n63_o;
  wire [2:0] n64_o;
  wire n65_o;
  wire n66_o;
  wire [12:0] n68_o;
  wire [6:0] n69_o;
  wire [5:0] n70_o;
  wire [3:0] n72_o;
  wire [4:0] n73_o;
  wire n74_o;
  wire [5:0] n75_o;
  wire [6:0] n77_o;
  wire [6:0] n78_o;
  wire [6:0] n79_o;
  wire [6:0] n80_o;
  wire [5:0] n81_o;
  wire [11:0] n82_o;
  wire [3:0] n83_o;
  wire n84_o;
  wire n85_o;
  wire [12:0] n87_o;
  wire [7:0] n88_o;
  wire [4:0] n89_o;
  wire [4:0] n91_o;
  wire [5:0] n92_o;
  wire n93_o;
  wire [6:0] n94_o;
  wire [7:0] n96_o;
  wire [7:0] n97_o;
  wire [7:0] n98_o;
  wire [7:0] n99_o;
  wire [6:0] n100_o;
  wire [11:0] n101_o;
  wire [4:0] n102_o;
  wire n103_o;
  wire n104_o;
  wire [12:0] n106_o;
  wire [8:0] n107_o;
  wire [3:0] n108_o;
  wire [5:0] n110_o;
  wire [6:0] n111_o;
  wire n112_o;
  wire [7:0] n113_o;
  wire [8:0] n115_o;
  wire [8:0] n116_o;
  wire [8:0] n117_o;
  wire [8:0] n118_o;
  wire [7:0] n119_o;
  wire [11:0] n120_o;
  wire [5:0] n121_o;
  wire n122_o;
  wire n123_o;
  wire [12:0] n125_o;
  wire [9:0] n126_o;
  wire [2:0] n127_o;
  wire [6:0] n129_o;
  wire [7:0] n130_o;
  wire n131_o;
  wire [8:0] n132_o;
  wire [9:0] n134_o;
  wire [9:0] n135_o;
  wire [9:0] n136_o;
  wire [9:0] n137_o;
  wire [8:0] n138_o;
  wire [11:0] n139_o;
  wire [6:0] n140_o;
  wire n141_o;
  wire n142_o;
  wire [12:0] n144_o;
  wire [10:0] n145_o;
  wire [1:0] n146_o;
  wire [7:0] n148_o;
  wire [8:0] n149_o;
  wire n150_o;
  wire [9:0] n151_o;
  wire [10:0] n153_o;
  wire [10:0] n154_o;
  wire [10:0] n155_o;
  wire [10:0] n156_o;
  wire [9:0] n157_o;
  wire [11:0] n158_o;
  wire [7:0] n159_o;
  wire n160_o;
  wire n161_o;
  wire [12:0] n163_o;
  wire [11:0] n164_o;
  wire n165_o;
  wire [8:0] n167_o;
  wire [9:0] n168_o;
  wire n169_o;
  wire [10:0] n170_o;
  wire [11:0] n172_o;
  wire [11:0] n173_o;
  wire [11:0] n174_o;
  wire [11:0] n175_o;
  wire [10:0] n176_o;
  wire [11:0] n177_o;
  wire [8:0] n178_o;
  wire n179_o;
  wire n180_o;
  wire [12:0] n182_o;
  wire [9:0] n184_o;
  wire [10:0] n185_o;
  wire n186_o;
  wire [11:0] n187_o;
  wire [12:0] n189_o;
  wire [12:0] n190_o;
  wire [12:0] n191_o;
  wire [12:0] n192_o;
  wire [11:0] n193_o;
  wire [9:0] n194_o;
  wire n195_o;
  wire n196_o;
  wire [10:0] n197_o;
  wire [7:0] n198_o;
  wire n199_o;
  wire [7:0] n201_o;
  wire [7:0] n202_o;
  wire [15:0] n203_o;
  wire n206_o;
  wire n209_o;
  wire n212_o;
  wire n215_o;
  wire [3:0] n217_o;
  reg [2:0] n218_o;
  wire [18:0] n219_o;
  reg [7:0] n220_q;
  reg [7:0] n221_q;
  reg n222_q;
  reg [7:0] n223_q;
  reg [4:0] n224_q;
  reg [7:0] n225_q;
  reg [4:0] n226_q;
  reg n227_q;
  reg [11:0] n228_q;
  reg n229_q;
  reg [11:0] n230_q;
  reg [8:0] n231_q;
  reg [2:0] n232_q;
  reg [2:0] n233_q;
  assign R = n219_o;
  assign fracx = n19_o; // (signal)
  assign ern0 = n22_o; // (signal)
  assign xsx = n23_o; // (signal)
  assign ern1 = n28_o; // (signal)
  assign ern1_d1 = n220_q; // (signal)
  assign ern1_d2 = n221_q; // (signal)
  assign fracxnorm = n35_o; // (signal)
  assign s0 = 2'b01; // (signal)
  assign t1 = n45_o; // (signal)
  assign d1 = n47_o; // (signal)
  assign t1s = n49_o; // (signal)
  assign t1s_h = n50_o; // (signal)
  assign t1s_l = n51_o; // (signal)
  assign u1 = n58_o; // (signal)
  assign t3_h = n60_o; // (signal)
  assign t2 = n63_o; // (signal)
  assign s1 = n64_o; // (signal)
  assign d2 = n66_o; // (signal)
  assign t2s = n68_o; // (signal)
  assign t2s_h = n69_o; // (signal)
  assign t2s_l = n70_o; // (signal)
  assign u2 = n77_o; // (signal)
  assign t4_h = n79_o; // (signal)
  assign t3 = n82_o; // (signal)
  assign s2 = n83_o; // (signal)
  assign d3 = n85_o; // (signal)
  assign d3_d1 = n222_q; // (signal)
  assign t3s = n87_o; // (signal)
  assign t3s_h = n88_o; // (signal)
  assign t3s_h_d1 = n223_q; // (signal)
  assign t3s_l = n89_o; // (signal)
  assign t3s_l_d1 = n224_q; // (signal)
  assign u3 = n96_o; // (signal)
  assign u3_d1 = n225_q; // (signal)
  assign t5_h = n98_o; // (signal)
  assign t4 = n101_o; // (signal)
  assign s3 = n102_o; // (signal)
  assign s3_d1 = n226_q; // (signal)
  assign d4 = n104_o; // (signal)
  assign t4s = n106_o; // (signal)
  assign t4s_h = n107_o; // (signal)
  assign t4s_l = n108_o; // (signal)
  assign u4 = n115_o; // (signal)
  assign t6_h = n117_o; // (signal)
  assign t5 = n120_o; // (signal)
  assign s4 = n121_o; // (signal)
  assign d5 = n123_o; // (signal)
  assign t5s = n125_o; // (signal)
  assign t5s_h = n126_o; // (signal)
  assign t5s_l = n127_o; // (signal)
  assign u5 = n134_o; // (signal)
  assign t7_h = n136_o; // (signal)
  assign t6 = n139_o; // (signal)
  assign s5 = n140_o; // (signal)
  assign d6 = n142_o; // (signal)
  assign t6s = n144_o; // (signal)
  assign t6s_h = n145_o; // (signal)
  assign t6s_l = n146_o; // (signal)
  assign u6 = n153_o; // (signal)
  assign t8_h = n155_o; // (signal)
  assign t7 = n158_o; // (signal)
  assign s6 = n159_o; // (signal)
  assign d7 = n161_o; // (signal)
  assign d7_d1 = n227_q; // (signal)
  assign t7s = n163_o; // (signal)
  assign t7s_h = n164_o; // (signal)
  assign t7s_h_d1 = n228_q; // (signal)
  assign t7s_l = n165_o; // (signal)
  assign t7s_l_d1 = n229_q; // (signal)
  assign u7 = n172_o; // (signal)
  assign u7_d1 = n230_q; // (signal)
  assign t9_h = n174_o; // (signal)
  assign t8 = n177_o; // (signal)
  assign s7 = n178_o; // (signal)
  assign s7_d1 = n231_q; // (signal)
  assign d8 = n180_o; // (signal)
  assign t8s = n182_o; // (signal)
  assign t8s_h = t8s; // (signal)
  assign u8 = n189_o; // (signal)
  assign t10_h = n191_o; // (signal)
  assign t9 = n193_o; // (signal)
  assign s8 = n194_o; // (signal)
  assign d10 = n196_o; // (signal)
  assign mr = n197_o; // (signal)
  assign fr = n198_o; // (signal)
  assign round = n199_o; // (signal)
  assign frrnd = n202_o; // (signal)
  assign rn2 = n203_o; // (signal)
  assign xsr = n218_o; // (signal)
  assign xsr_d1 = n232_q; // (signal)
  assign xsr_d2 = n233_q; // (signal)
  assign n19_o = X[7:0];
  assign n20_o = X[15:9];
  assign n22_o = {1'b0, n20_o};
  assign n23_o = X[18:16];
  assign n25_o = ern0 + 8'b00111111;
  assign n26_o = X[8];
  assign n27_o = {7'b0, n26_o};  //  uext
  assign n28_o = n25_o + n27_o;
  assign n30_o = {1'b1, fracx};
  assign n32_o = {n30_o, 3'b000};
  assign n33_o = X[8];
  assign n34_o = ~n33_o;
  assign n35_o = n34_o ? n32_o : n39_o;
  assign n37_o = {2'b01, fracx};
  assign n39_o = {n37_o, 2'b00};
  assign n41_o = fracxnorm[11:8];
  assign n43_o = 4'b0111 + n41_o;
  assign n44_o = fracxnorm[7:0];
  assign n45_o = {n43_o, n44_o};
  assign n46_o = t1[11];
  assign n47_o = ~n46_o;
  assign n49_o = {t1, 1'b0};
  assign n50_o = t1s[12:7];
  assign n51_o = t1s[6:0];
  assign n53_o = {1'b0, s0};
  assign n54_o = {n53_o, d1};
  assign n55_o = ~d1;
  assign n56_o = {n54_o, n55_o};
  assign n58_o = {n56_o, 1'b1};
  assign n59_o = t1s_h - u1;
  assign n60_o = d1 ? n59_o : n61_o;
  assign n61_o = t1s_h + u1;
  assign n62_o = t3_h[4:0];
  assign n63_o = {n62_o, t1s_l};
  assign n64_o = {s0, d1};
  assign n65_o = t2[11];
  assign n66_o = ~n65_o;
  assign n68_o = {t2, 1'b0};
  assign n69_o = t2s[12:6];
  assign n70_o = t2s[5:0];
  assign n72_o = {1'b0, s1};
  assign n73_o = {n72_o, d2};
  assign n74_o = ~d2;
  assign n75_o = {n73_o, n74_o};
  assign n77_o = {n75_o, 1'b1};
  assign n78_o = t2s_h - u2;
  assign n79_o = d2 ? n78_o : n80_o;
  assign n80_o = t2s_h + u2;
  assign n81_o = t4_h[5:0];
  assign n82_o = {n81_o, t2s_l};
  assign n83_o = {s1, d2};
  assign n84_o = t3[11];
  assign n85_o = ~n84_o;
  assign n87_o = {t3, 1'b0};
  assign n88_o = t3s[12:5];
  assign n89_o = t3s[4:0];
  assign n91_o = {1'b0, s2};
  assign n92_o = {n91_o, d3};
  assign n93_o = ~d3;
  assign n94_o = {n92_o, n93_o};
  assign n96_o = {n94_o, 1'b1};
  assign n97_o = t3s_h_d1 - u3_d1;
  assign n98_o = d3_d1 ? n97_o : n99_o;
  assign n99_o = t3s_h_d1 + u3_d1;
  assign n100_o = t5_h[6:0];
  assign n101_o = {n100_o, t3s_l_d1};
  assign n102_o = {s2, d3};
  assign n103_o = t4[11];
  assign n104_o = ~n103_o;
  assign n106_o = {t4, 1'b0};
  assign n107_o = t4s[12:4];
  assign n108_o = t4s[3:0];
  assign n110_o = {1'b0, s3_d1};
  assign n111_o = {n110_o, d4};
  assign n112_o = ~d4;
  assign n113_o = {n111_o, n112_o};
  assign n115_o = {n113_o, 1'b1};
  assign n116_o = t4s_h - u4;
  assign n117_o = d4 ? n116_o : n118_o;
  assign n118_o = t4s_h + u4;
  assign n119_o = t6_h[7:0];
  assign n120_o = {n119_o, t4s_l};
  assign n121_o = {s3_d1, d4};
  assign n122_o = t5[11];
  assign n123_o = ~n122_o;
  assign n125_o = {t5, 1'b0};
  assign n126_o = t5s[12:3];
  assign n127_o = t5s[2:0];
  assign n129_o = {1'b0, s4};
  assign n130_o = {n129_o, d5};
  assign n131_o = ~d5;
  assign n132_o = {n130_o, n131_o};
  assign n134_o = {n132_o, 1'b1};
  assign n135_o = t5s_h - u5;
  assign n136_o = d5 ? n135_o : n137_o;
  assign n137_o = t5s_h + u5;
  assign n138_o = t7_h[8:0];
  assign n139_o = {n138_o, t5s_l};
  assign n140_o = {s4, d5};
  assign n141_o = t6[11];
  assign n142_o = ~n141_o;
  assign n144_o = {t6, 1'b0};
  assign n145_o = t6s[12:2];
  assign n146_o = t6s[1:0];
  assign n148_o = {1'b0, s5};
  assign n149_o = {n148_o, d6};
  assign n150_o = ~d6;
  assign n151_o = {n149_o, n150_o};
  assign n153_o = {n151_o, 1'b1};
  assign n154_o = t6s_h - u6;
  assign n155_o = d6 ? n154_o : n156_o;
  assign n156_o = t6s_h + u6;
  assign n157_o = t8_h[9:0];
  assign n158_o = {n157_o, t6s_l};
  assign n159_o = {s5, d6};
  assign n160_o = t7[11];
  assign n161_o = ~n160_o;
  assign n163_o = {t7, 1'b0};
  assign n164_o = t7s[12:1];
  assign n165_o = t7s[0];
  assign n167_o = {1'b0, s6};
  assign n168_o = {n167_o, d7};
  assign n169_o = ~d7;
  assign n170_o = {n168_o, n169_o};
  assign n172_o = {n170_o, 1'b1};
  assign n173_o = t7s_h_d1 - u7_d1;
  assign n174_o = d7_d1 ? n173_o : n175_o;
  assign n175_o = t7s_h_d1 + u7_d1;
  assign n176_o = t9_h[10:0];
  assign n177_o = {n176_o, t7s_l_d1};
  assign n178_o = {s6, d7};
  assign n179_o = t8[11];
  assign n180_o = ~n179_o;
  assign n182_o = {t8, 1'b0};
  assign n184_o = {1'b0, s7_d1};
  assign n185_o = {n184_o, d8};
  assign n186_o = ~d8;
  assign n187_o = {n185_o, n186_o};
  assign n189_o = {n187_o, 1'b1};
  assign n190_o = t8s_h - u8;
  assign n191_o = d8 ? n190_o : n192_o;
  assign n192_o = t8s_h + u8;
  assign n193_o = t10_h[11:0];
  assign n194_o = {s7_d1, d8};
  assign n195_o = t9[11];
  assign n196_o = ~n195_o;
  assign n197_o = {s8, d10};
  assign n198_o = mr[8:1];
  assign n199_o = mr[0];
  assign n201_o = {7'b0000000, round};
  assign n202_o = fr + n201_o;
  assign n203_o = {ern1_d2, frrnd};
  assign n206_o = xsx == 3'b010;
  assign n209_o = xsx == 3'b100;
  assign n212_o = xsx == 3'b000;
  assign n215_o = xsx == 3'b001;
  assign n217_o = {n215_o, n212_o, n209_o, n206_o};
  always @*
    case (n217_o)
      4'b1000: n218_o = 3'b001;
      4'b0100: n218_o = 3'b000;
      4'b0010: n218_o = 3'b100;
      4'b0001: n218_o = 3'b010;
      default: n218_o = 3'b110;
    endcase
  assign n219_o = {xsr_d2, rn2};
  always @(posedge clk)
    n220_q <= ern1;
  always @(posedge clk)
    n221_q <= ern1_d1;
  always @(posedge clk)
    n222_q <= d3;
  always @(posedge clk)
    n223_q <= t3s_h;
  always @(posedge clk)
    n224_q <= t3s_l;
  always @(posedge clk)
    n225_q <= u3;
  always @(posedge clk)
    n226_q <= s3;
  always @(posedge clk)
    n227_q <= d7;
  always @(posedge clk)
    n228_q <= t7s_h;
  always @(posedge clk)
    n229_q <= t7s_l;
  always @(posedge clk)
    n230_q <= u7;
  always @(posedge clk)
    n231_q <= s7;
  always @(posedge clk)
    n232_q <= xsr;
  always @(posedge clk)
    n233_q <= xsr_d1;
endmodule

