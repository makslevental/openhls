module selfunction_f300_uid4
    (input wire[8:0] x,
        output wire[2:0] y);
    wire[2:0] y0;
    wire[2:0] y1;
    wire n303_o;
    wire n306_o;
    wire n309_o;
    wire n312_o;
    wire n315_o;
    wire n318_o;
    wire n321_o;
    wire n324_o;
    wire n327_o;
    wire n330_o;
    wire n333_o;
    wire n336_o;
    wire n339_o;
    wire n342_o;
    wire n345_o;
    wire n348_o;
    wire n351_o;
    wire n354_o;
    wire n357_o;
    wire n360_o;
    wire n363_o;
    wire n366_o;
    wire n369_o;
    wire n372_o;
    wire n375_o;
    wire n378_o;
    wire n381_o;
    wire n384_o;
    wire n387_o;
    wire n390_o;
    wire n393_o;
    wire n396_o;
    wire n399_o;
    wire n402_o;
    wire n405_o;
    wire n408_o;
    wire n411_o;
    wire n414_o;
    wire n417_o;
    wire n420_o;
    wire n423_o;
    wire n426_o;
    wire n429_o;
    wire n432_o;
    wire n435_o;
    wire n438_o;
    wire n441_o;
    wire n444_o;
    wire n447_o;
    wire n450_o;
    wire n453_o;
    wire n456_o;
    wire n459_o;
    wire n462_o;
    wire n465_o;
    wire n468_o;
    wire n471_o;
    wire n474_o;
    wire n477_o;
    wire n480_o;
    wire n483_o;
    wire n486_o;
    wire n489_o;
    wire n492_o;
    wire n495_o;
    wire n498_o;
    wire n501_o;
    wire n504_o;
    wire n507_o;
    wire n510_o;
    wire n513_o;
    wire n516_o;
    wire n519_o;
    wire n522_o;
    wire n525_o;
    wire n528_o;
    wire n531_o;
    wire n534_o;
    wire n537_o;
    wire n540_o;
    wire n543_o;
    wire n546_o;
    wire n549_o;
    wire n552_o;
    wire n555_o;
    wire n558_o;
    wire n561_o;
    wire n564_o;
    wire n567_o;
    wire n570_o;
    wire n573_o;
    wire n576_o;
    wire n579_o;
    wire n582_o;
    wire n585_o;
    wire n588_o;
    wire n591_o;
    wire n594_o;
    wire n597_o;
    wire n600_o;
    wire n603_o;
    wire n606_o;
    wire n609_o;
    wire n612_o;
    wire n615_o;
    wire n618_o;
    wire n621_o;
    wire n624_o;
    wire n627_o;
    wire n630_o;
    wire n633_o;
    wire n636_o;
    wire n639_o;
    wire n642_o;
    wire n645_o;
    wire n648_o;
    wire n651_o;
    wire n654_o;
    wire n657_o;
    wire n660_o;
    wire n663_o;
    wire n666_o;
    wire n669_o;
    wire n672_o;
    wire n675_o;
    wire n678_o;
    wire n681_o;
    wire n684_o;
    wire n687_o;
    wire n690_o;
    wire n693_o;
    wire n696_o;
    wire n699_o;
    wire n702_o;
    wire n705_o;
    wire n708_o;
    wire n711_o;
    wire n714_o;
    wire n717_o;
    wire n720_o;
    wire n723_o;
    wire n726_o;
    wire n729_o;
    wire n732_o;
    wire n735_o;
    wire n738_o;
    wire n741_o;
    wire n744_o;
    wire n747_o;
    wire n750_o;
    wire n753_o;
    wire n756_o;
    wire n759_o;
    wire n762_o;
    wire n765_o;
    wire n768_o;
    wire n771_o;
    wire n774_o;
    wire n777_o;
    wire n780_o;
    wire n783_o;
    wire n786_o;
    wire n789_o;
    wire n792_o;
    wire n795_o;
    wire n798_o;
    wire n801_o;
    wire n804_o;
    wire n807_o;
    wire n810_o;
    wire n813_o;
    wire n816_o;
    wire n819_o;
    wire n822_o;
    wire n825_o;
    wire n828_o;
    wire n831_o;
    wire n834_o;
    wire n837_o;
    wire n840_o;
    wire n843_o;
    wire n846_o;
    wire n849_o;
    wire n852_o;
    wire n855_o;
    wire n858_o;
    wire n861_o;
    wire n864_o;
    wire n867_o;
    wire n870_o;
    wire n873_o;
    wire n876_o;
    wire n879_o;
    wire n882_o;
    wire n885_o;
    wire n888_o;
    wire n891_o;
    wire n894_o;
    wire n897_o;
    wire n900_o;
    wire n903_o;
    wire n906_o;
    wire n909_o;
    wire n912_o;
    wire n915_o;
    wire n918_o;
    wire n921_o;
    wire n924_o;
    wire n927_o;
    wire n930_o;
    wire n933_o;
    wire n936_o;
    wire n939_o;
    wire n942_o;
    wire n945_o;
    wire n948_o;
    wire n951_o;
    wire n954_o;
    wire n957_o;
    wire n960_o;
    wire n963_o;
    wire n966_o;
    wire n969_o;
    wire n972_o;
    wire n975_o;
    wire n978_o;
    wire n981_o;
    wire n984_o;
    wire n987_o;
    wire n990_o;
    wire n993_o;
    wire n996_o;
    wire n999_o;
    wire n1002_o;
    wire n1005_o;
    wire n1008_o;
    wire n1011_o;
    wire n1014_o;
    wire n1017_o;
    wire n1020_o;
    wire n1023_o;
    wire n1026_o;
    wire n1029_o;
    wire n1032_o;
    wire n1035_o;
    wire n1038_o;
    wire n1041_o;
    wire n1044_o;
    wire n1047_o;
    wire n1050_o;
    wire n1053_o;
    wire n1056_o;
    wire n1059_o;
    wire n1062_o;
    wire n1065_o;
    wire n1068_o;
    wire n1071_o;
    wire n1074_o;
    wire n1077_o;
    wire n1080_o;
    wire n1083_o;
    wire n1086_o;
    wire n1089_o;
    wire n1092_o;
    wire n1095_o;
    wire n1098_o;
    wire n1101_o;
    wire n1104_o;
    wire n1107_o;
    wire n1110_o;
    wire n1113_o;
    wire n1116_o;
    wire n1119_o;
    wire n1122_o;
    wire n1125_o;
    wire n1128_o;
    wire n1131_o;
    wire n1134_o;
    wire n1137_o;
    wire n1140_o;
    wire n1143_o;
    wire n1146_o;
    wire n1149_o;
    wire n1152_o;
    wire n1155_o;
    wire n1158_o;
    wire n1161_o;
    wire n1164_o;
    wire n1167_o;
    wire n1170_o;
    wire n1173_o;
    wire n1176_o;
    wire n1179_o;
    wire n1182_o;
    wire n1185_o;
    wire n1188_o;
    wire n1191_o;
    wire n1194_o;
    wire n1197_o;
    wire n1200_o;
    wire n1203_o;
    wire n1206_o;
    wire n1209_o;
    wire n1212_o;
    wire n1215_o;
    wire n1218_o;
    wire n1221_o;
    wire n1224_o;
    wire n1227_o;
    wire n1230_o;
    wire n1233_o;
    wire n1236_o;
    wire n1239_o;
    wire n1242_o;
    wire n1245_o;
    wire n1248_o;
    wire n1251_o;
    wire n1254_o;
    wire n1257_o;
    wire n1260_o;
    wire n1263_o;
    wire n1266_o;
    wire n1269_o;
    wire n1272_o;
    wire n1275_o;
    wire n1278_o;
    wire n1281_o;
    wire n1284_o;
    wire n1287_o;
    wire n1290_o;
    wire n1293_o;
    wire n1296_o;
    wire n1299_o;
    wire n1302_o;
    wire n1305_o;
    wire n1308_o;
    wire n1311_o;
    wire n1314_o;
    wire n1317_o;
    wire n1320_o;
    wire n1323_o;
    wire n1326_o;
    wire n1329_o;
    wire n1332_o;
    wire n1335_o;
    wire n1338_o;
    wire n1341_o;
    wire n1344_o;
    wire n1347_o;
    wire n1350_o;
    wire n1353_o;
    wire n1356_o;
    wire n1359_o;
    wire n1362_o;
    wire n1365_o;
    wire n1368_o;
    wire n1371_o;
    wire n1374_o;
    wire n1377_o;
    wire n1380_o;
    wire n1383_o;
    wire n1386_o;
    wire n1389_o;
    wire n1392_o;
    wire n1395_o;
    wire n1398_o;
    wire n1401_o;
    wire n1404_o;
    wire n1407_o;
    wire n1410_o;
    wire n1413_o;
    wire n1416_o;
    wire n1419_o;
    wire n1422_o;
    wire n1425_o;
    wire n1428_o;
    wire n1431_o;
    wire n1434_o;
    wire n1437_o;
    wire n1440_o;
    wire n1443_o;
    wire n1446_o;
    wire n1449_o;
    wire n1452_o;
    wire n1455_o;
    wire n1458_o;
    wire n1461_o;
    wire n1464_o;
    wire n1467_o;
    wire n1470_o;
    wire n1473_o;
    wire n1476_o;
    wire n1479_o;
    wire n1482_o;
    wire n1485_o;
    wire n1488_o;
    wire n1491_o;
    wire n1494_o;
    wire n1497_o;
    wire n1500_o;
    wire n1503_o;
    wire n1506_o;
    wire n1509_o;
    wire n1512_o;
    wire n1515_o;
    wire n1518_o;
    wire n1521_o;
    wire n1524_o;
    wire n1527_o;
    wire n1530_o;
    wire n1533_o;
    wire n1536_o;
    wire n1539_o;
    wire n1542_o;
    wire n1545_o;
    wire n1548_o;
    wire n1551_o;
    wire n1554_o;
    wire n1557_o;
    wire n1560_o;
    wire n1563_o;
    wire n1566_o;
    wire n1569_o;
    wire n1572_o;
    wire n1575_o;
    wire n1578_o;
    wire n1581_o;
    wire n1584_o;
    wire n1587_o;
    wire n1590_o;
    wire n1593_o;
    wire n1596_o;
    wire n1599_o;
    wire n1602_o;
    wire n1605_o;
    wire n1608_o;
    wire n1611_o;
    wire n1614_o;
    wire n1617_o;
    wire n1620_o;
    wire n1623_o;
    wire n1626_o;
    wire n1629_o;
    wire n1632_o;
    wire n1635_o;
    wire n1638_o;
    wire n1641_o;
    wire n1644_o;
    wire n1647_o;
    wire n1650_o;
    wire n1653_o;
    wire n1656_o;
    wire n1659_o;
    wire n1662_o;
    wire n1665_o;
    wire n1668_o;
    wire n1671_o;
    wire n1674_o;
    wire n1677_o;
    wire n1680_o;
    wire n1683_o;
    wire n1686_o;
    wire n1689_o;
    wire n1692_o;
    wire n1695_o;
    wire n1698_o;
    wire n1701_o;
    wire n1704_o;
    wire n1707_o;
    wire n1710_o;
    wire n1713_o;
    wire n1716_o;
    wire n1719_o;
    wire n1722_o;
    wire n1725_o;
    wire n1728_o;
    wire n1731_o;
    wire n1734_o;
    wire n1737_o;
    wire n1740_o;
    wire n1743_o;
    wire n1746_o;
    wire n1749_o;
    wire n1752_o;
    wire n1755_o;
    wire n1758_o;
    wire n1761_o;
    wire n1764_o;
    wire n1767_o;
    wire n1770_o;
    wire n1773_o;
    wire n1776_o;
    wire n1779_o;
    wire n1782_o;
    wire n1785_o;
    wire n1788_o;
    wire n1791_o;
    wire n1794_o;
    wire n1797_o;
    wire n1800_o;
    wire n1803_o;
    wire n1806_o;
    wire n1809_o;
    wire n1812_o;
    wire n1815_o;
    wire n1818_o;
    wire n1821_o;
    wire n1824_o;
    wire n1827_o;
    wire n1830_o;
    wire n1833_o;
    wire n1836_o;
    wire[511:0] n1838_o;
    reg[2:0] n1839_o;
    assign y = y1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:28:8  */
    assign y0 = n1839_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:33:8  */
    assign y1 = y0; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:36:13  */
    assign n303_o = x == 9'b000000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:37:13  */
    assign n306_o = x == 9'b000000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:38:13  */
    assign n309_o = x == 9'b000000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:39:13  */
    assign n312_o = x == 9'b000000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:40:13  */
    assign n315_o = x == 9'b000000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:41:13  */
    assign n318_o = x == 9'b000000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:42:13  */
    assign n321_o = x == 9'b000000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:43:13  */
    assign n324_o = x == 9'b000000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:44:13  */
    assign n327_o = x == 9'b000001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:45:13  */
    assign n330_o = x == 9'b000001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:46:13  */
    assign n333_o = x == 9'b000001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:47:13  */
    assign n336_o = x == 9'b000001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:48:13  */
    assign n339_o = x == 9'b000001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:49:13  */
    assign n342_o = x == 9'b000001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:50:13  */
    assign n345_o = x == 9'b000001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:51:13  */
    assign n348_o = x == 9'b000001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:52:13  */
    assign n351_o = x == 9'b000010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:53:13  */
    assign n354_o = x == 9'b000010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:54:13  */
    assign n357_o = x == 9'b000010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:55:13  */
    assign n360_o = x == 9'b000010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:56:13  */
    assign n363_o = x == 9'b000010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:57:13  */
    assign n366_o = x == 9'b000010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:58:13  */
    assign n369_o = x == 9'b000010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:59:13  */
    assign n372_o = x == 9'b000010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:60:13  */
    assign n375_o = x == 9'b000011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:61:13  */
    assign n378_o = x == 9'b000011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:62:13  */
    assign n381_o = x == 9'b000011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:63:13  */
    assign n384_o = x == 9'b000011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:64:13  */
    assign n387_o = x == 9'b000011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:65:13  */
    assign n390_o = x == 9'b000011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:66:13  */
    assign n393_o = x == 9'b000011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:67:13  */
    assign n396_o = x == 9'b000011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:68:13  */
    assign n399_o = x == 9'b000100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:69:13  */
    assign n402_o = x == 9'b000100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:70:13  */
    assign n405_o = x == 9'b000100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:71:13  */
    assign n408_o = x == 9'b000100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:72:13  */
    assign n411_o = x == 9'b000100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:73:13  */
    assign n414_o = x == 9'b000100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:74:13  */
    assign n417_o = x == 9'b000100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:75:13  */
    assign n420_o = x == 9'b000100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:76:13  */
    assign n423_o = x == 9'b000101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:77:13  */
    assign n426_o = x == 9'b000101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:78:13  */
    assign n429_o = x == 9'b000101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:79:13  */
    assign n432_o = x == 9'b000101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:80:13  */
    assign n435_o = x == 9'b000101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:81:13  */
    assign n438_o = x == 9'b000101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:82:13  */
    assign n441_o = x == 9'b000101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:83:13  */
    assign n444_o = x == 9'b000101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:84:13  */
    assign n447_o = x == 9'b000110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:85:13  */
    assign n450_o = x == 9'b000110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:86:13  */
    assign n453_o = x == 9'b000110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:87:13  */
    assign n456_o = x == 9'b000110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:88:13  */
    assign n459_o = x == 9'b000110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:89:13  */
    assign n462_o = x == 9'b000110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:90:13  */
    assign n465_o = x == 9'b000110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:91:13  */
    assign n468_o = x == 9'b000110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:92:13  */
    assign n471_o = x == 9'b000111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:93:13  */
    assign n474_o = x == 9'b000111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:94:13  */
    assign n477_o = x == 9'b000111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:95:13  */
    assign n480_o = x == 9'b000111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:96:13  */
    assign n483_o = x == 9'b000111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:97:13  */
    assign n486_o = x == 9'b000111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:98:13  */
    assign n489_o = x == 9'b000111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:99:13  */
    assign n492_o = x == 9'b000111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:100:13  */
    assign n495_o = x == 9'b001000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:101:13  */
    assign n498_o = x == 9'b001000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:102:13  */
    assign n501_o = x == 9'b001000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:103:13  */
    assign n504_o = x == 9'b001000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:104:13  */
    assign n507_o = x == 9'b001000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:105:13  */
    assign n510_o = x == 9'b001000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:106:13  */
    assign n513_o = x == 9'b001000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:107:13  */
    assign n516_o = x == 9'b001000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:108:13  */
    assign n519_o = x == 9'b001001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:109:13  */
    assign n522_o = x == 9'b001001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:110:13  */
    assign n525_o = x == 9'b001001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:111:13  */
    assign n528_o = x == 9'b001001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:112:13  */
    assign n531_o = x == 9'b001001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:113:13  */
    assign n534_o = x == 9'b001001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:114:13  */
    assign n537_o = x == 9'b001001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:115:13  */
    assign n540_o = x == 9'b001001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:116:13  */
    assign n543_o = x == 9'b001010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:117:13  */
    assign n546_o = x == 9'b001010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:118:13  */
    assign n549_o = x == 9'b001010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:119:13  */
    assign n552_o = x == 9'b001010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:120:13  */
    assign n555_o = x == 9'b001010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:121:13  */
    assign n558_o = x == 9'b001010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:122:13  */
    assign n561_o = x == 9'b001010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:123:13  */
    assign n564_o = x == 9'b001010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:124:13  */
    assign n567_o = x == 9'b001011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:125:13  */
    assign n570_o = x == 9'b001011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:126:13  */
    assign n573_o = x == 9'b001011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:127:13  */
    assign n576_o = x == 9'b001011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:128:13  */
    assign n579_o = x == 9'b001011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:129:13  */
    assign n582_o = x == 9'b001011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:130:13  */
    assign n585_o = x == 9'b001011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:131:13  */
    assign n588_o = x == 9'b001011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:132:13  */
    assign n591_o = x == 9'b001100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:133:13  */
    assign n594_o = x == 9'b001100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:134:13  */
    assign n597_o = x == 9'b001100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:135:13  */
    assign n600_o = x == 9'b001100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:136:13  */
    assign n603_o = x == 9'b001100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:137:13  */
    assign n606_o = x == 9'b001100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:138:13  */
    assign n609_o = x == 9'b001100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:139:13  */
    assign n612_o = x == 9'b001100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:140:13  */
    assign n615_o = x == 9'b001101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:141:13  */
    assign n618_o = x == 9'b001101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:142:13  */
    assign n621_o = x == 9'b001101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:143:13  */
    assign n624_o = x == 9'b001101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:144:13  */
    assign n627_o = x == 9'b001101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:145:13  */
    assign n630_o = x == 9'b001101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:146:13  */
    assign n633_o = x == 9'b001101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:147:13  */
    assign n636_o = x == 9'b001101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:148:13  */
    assign n639_o = x == 9'b001110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:149:13  */
    assign n642_o = x == 9'b001110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:150:13  */
    assign n645_o = x == 9'b001110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:151:13  */
    assign n648_o = x == 9'b001110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:152:13  */
    assign n651_o = x == 9'b001110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:153:13  */
    assign n654_o = x == 9'b001110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:154:13  */
    assign n657_o = x == 9'b001110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:155:13  */
    assign n660_o = x == 9'b001110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:156:13  */
    assign n663_o = x == 9'b001111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:157:13  */
    assign n666_o = x == 9'b001111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:158:13  */
    assign n669_o = x == 9'b001111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:159:13  */
    assign n672_o = x == 9'b001111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:160:13  */
    assign n675_o = x == 9'b001111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:161:13  */
    assign n678_o = x == 9'b001111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:162:13  */
    assign n681_o = x == 9'b001111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:163:13  */
    assign n684_o = x == 9'b001111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:164:13  */
    assign n687_o = x == 9'b010000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:165:13  */
    assign n690_o = x == 9'b010000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:166:13  */
    assign n693_o = x == 9'b010000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:167:13  */
    assign n696_o = x == 9'b010000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:168:13  */
    assign n699_o = x == 9'b010000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:169:13  */
    assign n702_o = x == 9'b010000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:170:13  */
    assign n705_o = x == 9'b010000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:171:13  */
    assign n708_o = x == 9'b010000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:172:13  */
    assign n711_o = x == 9'b010001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:173:13  */
    assign n714_o = x == 9'b010001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:174:13  */
    assign n717_o = x == 9'b010001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:175:13  */
    assign n720_o = x == 9'b010001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:176:13  */
    assign n723_o = x == 9'b010001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:177:13  */
    assign n726_o = x == 9'b010001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:178:13  */
    assign n729_o = x == 9'b010001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:179:13  */
    assign n732_o = x == 9'b010001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:180:13  */
    assign n735_o = x == 9'b010010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:181:13  */
    assign n738_o = x == 9'b010010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:182:13  */
    assign n741_o = x == 9'b010010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:183:13  */
    assign n744_o = x == 9'b010010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:184:13  */
    assign n747_o = x == 9'b010010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:185:13  */
    assign n750_o = x == 9'b010010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:186:13  */
    assign n753_o = x == 9'b010010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:187:13  */
    assign n756_o = x == 9'b010010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:188:13  */
    assign n759_o = x == 9'b010011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:189:13  */
    assign n762_o = x == 9'b010011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:190:13  */
    assign n765_o = x == 9'b010011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:191:13  */
    assign n768_o = x == 9'b010011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:192:13  */
    assign n771_o = x == 9'b010011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:193:13  */
    assign n774_o = x == 9'b010011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:194:13  */
    assign n777_o = x == 9'b010011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:195:13  */
    assign n780_o = x == 9'b010011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:196:13  */
    assign n783_o = x == 9'b010100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:197:13  */
    assign n786_o = x == 9'b010100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:198:13  */
    assign n789_o = x == 9'b010100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:199:13  */
    assign n792_o = x == 9'b010100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:200:13  */
    assign n795_o = x == 9'b010100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:201:13  */
    assign n798_o = x == 9'b010100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:202:13  */
    assign n801_o = x == 9'b010100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:203:13  */
    assign n804_o = x == 9'b010100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:204:13  */
    assign n807_o = x == 9'b010101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:205:13  */
    assign n810_o = x == 9'b010101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:206:13  */
    assign n813_o = x == 9'b010101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:207:13  */
    assign n816_o = x == 9'b010101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:208:13  */
    assign n819_o = x == 9'b010101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:209:13  */
    assign n822_o = x == 9'b010101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:210:13  */
    assign n825_o = x == 9'b010101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:211:13  */
    assign n828_o = x == 9'b010101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:212:13  */
    assign n831_o = x == 9'b010110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:213:13  */
    assign n834_o = x == 9'b010110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:214:13  */
    assign n837_o = x == 9'b010110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:215:13  */
    assign n840_o = x == 9'b010110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:216:13  */
    assign n843_o = x == 9'b010110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:217:13  */
    assign n846_o = x == 9'b010110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:218:13  */
    assign n849_o = x == 9'b010110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:219:13  */
    assign n852_o = x == 9'b010110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:220:13  */
    assign n855_o = x == 9'b010111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:221:13  */
    assign n858_o = x == 9'b010111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:222:13  */
    assign n861_o = x == 9'b010111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:223:13  */
    assign n864_o = x == 9'b010111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:224:13  */
    assign n867_o = x == 9'b010111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:225:13  */
    assign n870_o = x == 9'b010111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:226:13  */
    assign n873_o = x == 9'b010111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:227:13  */
    assign n876_o = x == 9'b010111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:228:13  */
    assign n879_o = x == 9'b011000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:229:13  */
    assign n882_o = x == 9'b011000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:230:13  */
    assign n885_o = x == 9'b011000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:231:13  */
    assign n888_o = x == 9'b011000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:232:13  */
    assign n891_o = x == 9'b011000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:233:13  */
    assign n894_o = x == 9'b011000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:234:13  */
    assign n897_o = x == 9'b011000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:235:13  */
    assign n900_o = x == 9'b011000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:236:13  */
    assign n903_o = x == 9'b011001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:237:13  */
    assign n906_o = x == 9'b011001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:238:13  */
    assign n909_o = x == 9'b011001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:239:13  */
    assign n912_o = x == 9'b011001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:240:13  */
    assign n915_o = x == 9'b011001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:241:13  */
    assign n918_o = x == 9'b011001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:242:13  */
    assign n921_o = x == 9'b011001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:243:13  */
    assign n924_o = x == 9'b011001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:244:13  */
    assign n927_o = x == 9'b011010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:245:13  */
    assign n930_o = x == 9'b011010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:246:13  */
    assign n933_o = x == 9'b011010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:247:13  */
    assign n936_o = x == 9'b011010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:248:13  */
    assign n939_o = x == 9'b011010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:249:13  */
    assign n942_o = x == 9'b011010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:250:13  */
    assign n945_o = x == 9'b011010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:251:13  */
    assign n948_o = x == 9'b011010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:252:13  */
    assign n951_o = x == 9'b011011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:253:13  */
    assign n954_o = x == 9'b011011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:254:13  */
    assign n957_o = x == 9'b011011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:255:13  */
    assign n960_o = x == 9'b011011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:256:13  */
    assign n963_o = x == 9'b011011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:257:13  */
    assign n966_o = x == 9'b011011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:258:13  */
    assign n969_o = x == 9'b011011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:259:13  */
    assign n972_o = x == 9'b011011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:260:13  */
    assign n975_o = x == 9'b011100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:261:13  */
    assign n978_o = x == 9'b011100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:262:13  */
    assign n981_o = x == 9'b011100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:263:13  */
    assign n984_o = x == 9'b011100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:264:13  */
    assign n987_o = x == 9'b011100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:265:13  */
    assign n990_o = x == 9'b011100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:266:13  */
    assign n993_o = x == 9'b011100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:267:13  */
    assign n996_o = x == 9'b011100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:268:13  */
    assign n999_o = x == 9'b011101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:269:13  */
    assign n1002_o = x == 9'b011101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:270:13  */
    assign n1005_o = x == 9'b011101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:271:13  */
    assign n1008_o = x == 9'b011101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:272:13  */
    assign n1011_o = x == 9'b011101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:273:13  */
    assign n1014_o = x == 9'b011101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:274:13  */
    assign n1017_o = x == 9'b011101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:275:13  */
    assign n1020_o = x == 9'b011101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:276:13  */
    assign n1023_o = x == 9'b011110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:277:13  */
    assign n1026_o = x == 9'b011110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:278:13  */
    assign n1029_o = x == 9'b011110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:279:13  */
    assign n1032_o = x == 9'b011110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:280:13  */
    assign n1035_o = x == 9'b011110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:281:13  */
    assign n1038_o = x == 9'b011110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:282:13  */
    assign n1041_o = x == 9'b011110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:283:13  */
    assign n1044_o = x == 9'b011110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:284:13  */
    assign n1047_o = x == 9'b011111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:285:13  */
    assign n1050_o = x == 9'b011111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:286:13  */
    assign n1053_o = x == 9'b011111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:287:13  */
    assign n1056_o = x == 9'b011111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:288:13  */
    assign n1059_o = x == 9'b011111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:289:13  */
    assign n1062_o = x == 9'b011111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:290:13  */
    assign n1065_o = x == 9'b011111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:291:13  */
    assign n1068_o = x == 9'b011111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:292:13  */
    assign n1071_o = x == 9'b100000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:293:13  */
    assign n1074_o = x == 9'b100000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:294:13  */
    assign n1077_o = x == 9'b100000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:295:13  */
    assign n1080_o = x == 9'b100000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:296:13  */
    assign n1083_o = x == 9'b100000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:297:13  */
    assign n1086_o = x == 9'b100000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:298:13  */
    assign n1089_o = x == 9'b100000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:299:13  */
    assign n1092_o = x == 9'b100000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:300:13  */
    assign n1095_o = x == 9'b100001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:301:13  */
    assign n1098_o = x == 9'b100001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:302:13  */
    assign n1101_o = x == 9'b100001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:303:13  */
    assign n1104_o = x == 9'b100001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:304:13  */
    assign n1107_o = x == 9'b100001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:305:13  */
    assign n1110_o = x == 9'b100001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:306:13  */
    assign n1113_o = x == 9'b100001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:307:13  */
    assign n1116_o = x == 9'b100001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:308:13  */
    assign n1119_o = x == 9'b100010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:309:13  */
    assign n1122_o = x == 9'b100010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:310:13  */
    assign n1125_o = x == 9'b100010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:311:13  */
    assign n1128_o = x == 9'b100010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:312:13  */
    assign n1131_o = x == 9'b100010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:313:13  */
    assign n1134_o = x == 9'b100010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:314:13  */
    assign n1137_o = x == 9'b100010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:315:13  */
    assign n1140_o = x == 9'b100010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:316:13  */
    assign n1143_o = x == 9'b100011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:317:13  */
    assign n1146_o = x == 9'b100011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:318:13  */
    assign n1149_o = x == 9'b100011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:319:13  */
    assign n1152_o = x == 9'b100011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:320:13  */
    assign n1155_o = x == 9'b100011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:321:13  */
    assign n1158_o = x == 9'b100011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:322:13  */
    assign n1161_o = x == 9'b100011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:323:13  */
    assign n1164_o = x == 9'b100011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:324:13  */
    assign n1167_o = x == 9'b100100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:325:13  */
    assign n1170_o = x == 9'b100100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:326:13  */
    assign n1173_o = x == 9'b100100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:327:13  */
    assign n1176_o = x == 9'b100100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:328:13  */
    assign n1179_o = x == 9'b100100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:329:13  */
    assign n1182_o = x == 9'b100100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:330:13  */
    assign n1185_o = x == 9'b100100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:331:13  */
    assign n1188_o = x == 9'b100100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:332:13  */
    assign n1191_o = x == 9'b100101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:333:13  */
    assign n1194_o = x == 9'b100101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:334:13  */
    assign n1197_o = x == 9'b100101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:335:13  */
    assign n1200_o = x == 9'b100101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:336:13  */
    assign n1203_o = x == 9'b100101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:337:13  */
    assign n1206_o = x == 9'b100101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:338:13  */
    assign n1209_o = x == 9'b100101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:339:13  */
    assign n1212_o = x == 9'b100101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:340:13  */
    assign n1215_o = x == 9'b100110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:341:13  */
    assign n1218_o = x == 9'b100110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:342:13  */
    assign n1221_o = x == 9'b100110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:343:13  */
    assign n1224_o = x == 9'b100110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:344:13  */
    assign n1227_o = x == 9'b100110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:345:13  */
    assign n1230_o = x == 9'b100110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:346:13  */
    assign n1233_o = x == 9'b100110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:347:13  */
    assign n1236_o = x == 9'b100110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:348:13  */
    assign n1239_o = x == 9'b100111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:349:13  */
    assign n1242_o = x == 9'b100111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:350:13  */
    assign n1245_o = x == 9'b100111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:351:13  */
    assign n1248_o = x == 9'b100111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:352:13  */
    assign n1251_o = x == 9'b100111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:353:13  */
    assign n1254_o = x == 9'b100111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:354:13  */
    assign n1257_o = x == 9'b100111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:355:13  */
    assign n1260_o = x == 9'b100111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:356:13  */
    assign n1263_o = x == 9'b101000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:357:13  */
    assign n1266_o = x == 9'b101000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:358:13  */
    assign n1269_o = x == 9'b101000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:359:13  */
    assign n1272_o = x == 9'b101000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:360:13  */
    assign n1275_o = x == 9'b101000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:361:13  */
    assign n1278_o = x == 9'b101000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:362:13  */
    assign n1281_o = x == 9'b101000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:363:13  */
    assign n1284_o = x == 9'b101000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:364:13  */
    assign n1287_o = x == 9'b101001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:365:13  */
    assign n1290_o = x == 9'b101001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:366:13  */
    assign n1293_o = x == 9'b101001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:367:13  */
    assign n1296_o = x == 9'b101001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:368:13  */
    assign n1299_o = x == 9'b101001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:369:13  */
    assign n1302_o = x == 9'b101001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:370:13  */
    assign n1305_o = x == 9'b101001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:371:13  */
    assign n1308_o = x == 9'b101001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:372:13  */
    assign n1311_o = x == 9'b101010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:373:13  */
    assign n1314_o = x == 9'b101010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:374:13  */
    assign n1317_o = x == 9'b101010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:375:13  */
    assign n1320_o = x == 9'b101010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:376:13  */
    assign n1323_o = x == 9'b101010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:377:13  */
    assign n1326_o = x == 9'b101010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:378:13  */
    assign n1329_o = x == 9'b101010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:379:13  */
    assign n1332_o = x == 9'b101010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:380:13  */
    assign n1335_o = x == 9'b101011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:381:13  */
    assign n1338_o = x == 9'b101011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:382:13  */
    assign n1341_o = x == 9'b101011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:383:13  */
    assign n1344_o = x == 9'b101011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:384:13  */
    assign n1347_o = x == 9'b101011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:385:13  */
    assign n1350_o = x == 9'b101011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:386:13  */
    assign n1353_o = x == 9'b101011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:387:13  */
    assign n1356_o = x == 9'b101011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:388:13  */
    assign n1359_o = x == 9'b101100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:389:13  */
    assign n1362_o = x == 9'b101100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:390:13  */
    assign n1365_o = x == 9'b101100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:391:13  */
    assign n1368_o = x == 9'b101100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:392:13  */
    assign n1371_o = x == 9'b101100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:393:13  */
    assign n1374_o = x == 9'b101100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:394:13  */
    assign n1377_o = x == 9'b101100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:395:13  */
    assign n1380_o = x == 9'b101100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:396:13  */
    assign n1383_o = x == 9'b101101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:397:13  */
    assign n1386_o = x == 9'b101101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:398:13  */
    assign n1389_o = x == 9'b101101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:399:13  */
    assign n1392_o = x == 9'b101101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:400:13  */
    assign n1395_o = x == 9'b101101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:401:13  */
    assign n1398_o = x == 9'b101101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:402:13  */
    assign n1401_o = x == 9'b101101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:403:13  */
    assign n1404_o = x == 9'b101101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:404:13  */
    assign n1407_o = x == 9'b101110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:405:13  */
    assign n1410_o = x == 9'b101110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:406:13  */
    assign n1413_o = x == 9'b101110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:407:13  */
    assign n1416_o = x == 9'b101110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:408:13  */
    assign n1419_o = x == 9'b101110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:409:13  */
    assign n1422_o = x == 9'b101110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:410:13  */
    assign n1425_o = x == 9'b101110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:411:13  */
    assign n1428_o = x == 9'b101110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:412:13  */
    assign n1431_o = x == 9'b101111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:413:13  */
    assign n1434_o = x == 9'b101111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:414:13  */
    assign n1437_o = x == 9'b101111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:415:13  */
    assign n1440_o = x == 9'b101111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:416:13  */
    assign n1443_o = x == 9'b101111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:417:13  */
    assign n1446_o = x == 9'b101111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:418:13  */
    assign n1449_o = x == 9'b101111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:419:13  */
    assign n1452_o = x == 9'b101111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:420:13  */
    assign n1455_o = x == 9'b110000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:421:13  */
    assign n1458_o = x == 9'b110000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:422:13  */
    assign n1461_o = x == 9'b110000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:423:13  */
    assign n1464_o = x == 9'b110000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:424:13  */
    assign n1467_o = x == 9'b110000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:425:13  */
    assign n1470_o = x == 9'b110000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:426:13  */
    assign n1473_o = x == 9'b110000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:427:13  */
    assign n1476_o = x == 9'b110000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:428:13  */
    assign n1479_o = x == 9'b110001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:429:13  */
    assign n1482_o = x == 9'b110001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:430:13  */
    assign n1485_o = x == 9'b110001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:431:13  */
    assign n1488_o = x == 9'b110001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:432:13  */
    assign n1491_o = x == 9'b110001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:433:13  */
    assign n1494_o = x == 9'b110001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:434:13  */
    assign n1497_o = x == 9'b110001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:435:13  */
    assign n1500_o = x == 9'b110001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:436:13  */
    assign n1503_o = x == 9'b110010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:437:13  */
    assign n1506_o = x == 9'b110010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:438:13  */
    assign n1509_o = x == 9'b110010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:439:13  */
    assign n1512_o = x == 9'b110010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:440:13  */
    assign n1515_o = x == 9'b110010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:441:13  */
    assign n1518_o = x == 9'b110010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:442:13  */
    assign n1521_o = x == 9'b110010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:443:13  */
    assign n1524_o = x == 9'b110010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:444:13  */
    assign n1527_o = x == 9'b110011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:445:13  */
    assign n1530_o = x == 9'b110011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:446:13  */
    assign n1533_o = x == 9'b110011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:447:13  */
    assign n1536_o = x == 9'b110011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:448:13  */
    assign n1539_o = x == 9'b110011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:449:13  */
    assign n1542_o = x == 9'b110011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:450:13  */
    assign n1545_o = x == 9'b110011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:451:13  */
    assign n1548_o = x == 9'b110011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:452:13  */
    assign n1551_o = x == 9'b110100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:453:13  */
    assign n1554_o = x == 9'b110100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:454:13  */
    assign n1557_o = x == 9'b110100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:455:13  */
    assign n1560_o = x == 9'b110100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:456:13  */
    assign n1563_o = x == 9'b110100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:457:13  */
    assign n1566_o = x == 9'b110100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:458:13  */
    assign n1569_o = x == 9'b110100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:459:13  */
    assign n1572_o = x == 9'b110100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:460:13  */
    assign n1575_o = x == 9'b110101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:461:13  */
    assign n1578_o = x == 9'b110101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:462:13  */
    assign n1581_o = x == 9'b110101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:463:13  */
    assign n1584_o = x == 9'b110101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:464:13  */
    assign n1587_o = x == 9'b110101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:465:13  */
    assign n1590_o = x == 9'b110101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:466:13  */
    assign n1593_o = x == 9'b110101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:467:13  */
    assign n1596_o = x == 9'b110101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:468:13  */
    assign n1599_o = x == 9'b110110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:469:13  */
    assign n1602_o = x == 9'b110110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:470:13  */
    assign n1605_o = x == 9'b110110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:471:13  */
    assign n1608_o = x == 9'b110110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:472:13  */
    assign n1611_o = x == 9'b110110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:473:13  */
    assign n1614_o = x == 9'b110110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:474:13  */
    assign n1617_o = x == 9'b110110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:475:13  */
    assign n1620_o = x == 9'b110110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:476:13  */
    assign n1623_o = x == 9'b110111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:477:13  */
    assign n1626_o = x == 9'b110111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:478:13  */
    assign n1629_o = x == 9'b110111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:479:13  */
    assign n1632_o = x == 9'b110111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:480:13  */
    assign n1635_o = x == 9'b110111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:481:13  */
    assign n1638_o = x == 9'b110111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:482:13  */
    assign n1641_o = x == 9'b110111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:483:13  */
    assign n1644_o = x == 9'b110111111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:484:13  */
    assign n1647_o = x == 9'b111000000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:485:13  */
    assign n1650_o = x == 9'b111000001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:486:13  */
    assign n1653_o = x == 9'b111000010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:487:13  */
    assign n1656_o = x == 9'b111000011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:488:13  */
    assign n1659_o = x == 9'b111000100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:489:13  */
    assign n1662_o = x == 9'b111000101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:490:13  */
    assign n1665_o = x == 9'b111000110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:491:13  */
    assign n1668_o = x == 9'b111000111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:492:13  */
    assign n1671_o = x == 9'b111001000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:493:13  */
    assign n1674_o = x == 9'b111001001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:494:13  */
    assign n1677_o = x == 9'b111001010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:495:13  */
    assign n1680_o = x == 9'b111001011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:496:13  */
    assign n1683_o = x == 9'b111001100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:497:13  */
    assign n1686_o = x == 9'b111001101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:498:13  */
    assign n1689_o = x == 9'b111001110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:499:13  */
    assign n1692_o = x == 9'b111001111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:500:13  */
    assign n1695_o = x == 9'b111010000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:501:13  */
    assign n1698_o = x == 9'b111010001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:502:13  */
    assign n1701_o = x == 9'b111010010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:503:13  */
    assign n1704_o = x == 9'b111010011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:504:13  */
    assign n1707_o = x == 9'b111010100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:505:13  */
    assign n1710_o = x == 9'b111010101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:506:13  */
    assign n1713_o = x == 9'b111010110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:507:13  */
    assign n1716_o = x == 9'b111010111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:508:13  */
    assign n1719_o = x == 9'b111011000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:509:13  */
    assign n1722_o = x == 9'b111011001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:510:13  */
    assign n1725_o = x == 9'b111011010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:511:13  */
    assign n1728_o = x == 9'b111011011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:512:13  */
    assign n1731_o = x == 9'b111011100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:513:13  */
    assign n1734_o = x == 9'b111011101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:514:13  */
    assign n1737_o = x == 9'b111011110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:515:13  */
    assign n1740_o = x == 9'b111011111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:516:13  */
    assign n1743_o = x == 9'b111100000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:517:13  */
    assign n1746_o = x == 9'b111100001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:518:13  */
    assign n1749_o = x == 9'b111100010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:519:13  */
    assign n1752_o = x == 9'b111100011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:520:13  */
    assign n1755_o = x == 9'b111100100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:521:13  */
    assign n1758_o = x == 9'b111100101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:522:13  */
    assign n1761_o = x == 9'b111100110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:523:13  */
    assign n1764_o = x == 9'b111100111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:524:13  */
    assign n1767_o = x == 9'b111101000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:525:13  */
    assign n1770_o = x == 9'b111101001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:526:13  */
    assign n1773_o = x == 9'b111101010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:527:13  */
    assign n1776_o = x == 9'b111101011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:528:13  */
    assign n1779_o = x == 9'b111101100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:529:13  */
    assign n1782_o = x == 9'b111101101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:530:13  */
    assign n1785_o = x == 9'b111101110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:531:13  */
    assign n1788_o = x == 9'b111101111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:532:13  */
    assign n1791_o = x == 9'b111110000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:533:13  */
    assign n1794_o = x == 9'b111110001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:534:13  */
    assign n1797_o = x == 9'b111110010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:535:13  */
    assign n1800_o = x == 9'b111110011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:536:13  */
    assign n1803_o = x == 9'b111110100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:537:13  */
    assign n1806_o = x == 9'b111110101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:538:13  */
    assign n1809_o = x == 9'b111110110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:539:13  */
    assign n1812_o = x == 9'b111110111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:540:13  */
    assign n1815_o = x == 9'b111111000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:541:13  */
    assign n1818_o = x == 9'b111111001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:542:13  */
    assign n1821_o = x == 9'b111111010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:543:13  */
    assign n1824_o = x == 9'b111111011;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:544:13  */
    assign n1827_o = x == 9'b111111100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:545:13  */
    assign n1830_o = x == 9'b111111101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:546:13  */
    assign n1833_o = x == 9'b111111110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:547:13  */
    assign n1836_o = x == 9'b111111111;
    assign n1838_o = {n1836_o, n1833_o, n1830_o, n1827_o, n1824_o, n1821_o, n1818_o, n1815_o, n1812_o, n1809_o, n1806_o, n1803_o, n1800_o, n1797_o, n1794_o, n1791_o, n1788_o, n1785_o, n1782_o, n1779_o, n1776_o, n1773_o, n1770_o, n1767_o, n1764_o, n1761_o, n1758_o, n1755_o, n1752_o, n1749_o, n1746_o, n1743_o, n1740_o, n1737_o, n1734_o, n1731_o, n1728_o, n1725_o, n1722_o, n1719_o, n1716_o, n1713_o, n1710_o, n1707_o, n1704_o, n1701_o, n1698_o, n1695_o, n1692_o, n1689_o, n1686_o, n1683_o, n1680_o, n1677_o, n1674_o, n1671_o, n1668_o, n1665_o, n1662_o, n1659_o, n1656_o, n1653_o, n1650_o, n1647_o, n1644_o, n1641_o, n1638_o, n1635_o, n1632_o, n1629_o, n1626_o, n1623_o, n1620_o, n1617_o, n1614_o, n1611_o, n1608_o, n1605_o, n1602_o, n1599_o, n1596_o, n1593_o, n1590_o, n1587_o, n1584_o, n1581_o, n1578_o, n1575_o, n1572_o, n1569_o, n1566_o, n1563_o, n1560_o, n1557_o, n1554_o, n1551_o, n1548_o, n1545_o, n1542_o, n1539_o, n1536_o, n1533_o, n1530_o, n1527_o, n1524_o, n1521_o, n1518_o, n1515_o, n1512_o, n1509_o, n1506_o, n1503_o, n1500_o, n1497_o, n1494_o, n1491_o, n1488_o, n1485_o, n1482_o, n1479_o, n1476_o, n1473_o, n1470_o, n1467_o, n1464_o, n1461_o, n1458_o, n1455_o, n1452_o, n1449_o, n1446_o, n1443_o, n1440_o, n1437_o, n1434_o, n1431_o, n1428_o, n1425_o, n1422_o, n1419_o, n1416_o, n1413_o, n1410_o, n1407_o, n1404_o, n1401_o, n1398_o, n1395_o, n1392_o, n1389_o, n1386_o, n1383_o, n1380_o, n1377_o, n1374_o, n1371_o, n1368_o, n1365_o, n1362_o, n1359_o, n1356_o, n1353_o, n1350_o, n1347_o, n1344_o, n1341_o, n1338_o, n1335_o, n1332_o, n1329_o, n1326_o, n1323_o, n1320_o, n1317_o, n1314_o, n1311_o, n1308_o, n1305_o, n1302_o, n1299_o, n1296_o, n1293_o, n1290_o, n1287_o, n1284_o, n1281_o, n1278_o, n1275_o, n1272_o, n1269_o, n1266_o, n1263_o, n1260_o, n1257_o, n1254_o, n1251_o, n1248_o, n1245_o, n1242_o, n1239_o, n1236_o, n1233_o, n1230_o, n1227_o, n1224_o, n1221_o, n1218_o, n1215_o, n1212_o, n1209_o, n1206_o, n1203_o, n1200_o, n1197_o, n1194_o, n1191_o, n1188_o, n1185_o, n1182_o, n1179_o, n1176_o, n1173_o, n1170_o, n1167_o, n1164_o, n1161_o, n1158_o, n1155_o, n1152_o, n1149_o, n1146_o, n1143_o, n1140_o, n1137_o, n1134_o, n1131_o, n1128_o, n1125_o, n1122_o, n1119_o, n1116_o, n1113_o, n1110_o, n1107_o, n1104_o, n1101_o, n1098_o, n1095_o, n1092_o, n1089_o, n1086_o, n1083_o, n1080_o, n1077_o, n1074_o, n1071_o, n1068_o, n1065_o, n1062_o, n1059_o, n1056_o, n1053_o, n1050_o, n1047_o, n1044_o, n1041_o, n1038_o, n1035_o, n1032_o, n1029_o, n1026_o, n1023_o, n1020_o, n1017_o, n1014_o, n1011_o, n1008_o, n1005_o, n1002_o, n999_o, n996_o, n993_o, n990_o, n987_o, n984_o, n981_o, n978_o, n975_o, n972_o, n969_o, n966_o, n963_o, n960_o, n957_o, n954_o, n951_o, n948_o, n945_o, n942_o, n939_o, n936_o, n933_o, n930_o, n927_o, n924_o, n921_o, n918_o, n915_o, n912_o, n909_o, n906_o, n903_o, n900_o, n897_o, n894_o, n891_o, n888_o, n885_o, n882_o, n879_o, n876_o, n873_o, n870_o, n867_o, n864_o, n861_o, n858_o, n855_o, n852_o, n849_o, n846_o, n843_o, n840_o, n837_o, n834_o, n831_o, n828_o, n825_o, n822_o, n819_o, n816_o, n813_o, n810_o, n807_o, n804_o, n801_o, n798_o, n795_o, n792_o, n789_o, n786_o, n783_o, n780_o, n777_o, n774_o, n771_o, n768_o, n765_o, n762_o, n759_o, n756_o, n753_o, n750_o, n747_o, n744_o, n741_o, n738_o, n735_o, n732_o, n729_o, n726_o, n723_o, n720_o, n717_o, n714_o, n711_o, n708_o, n705_o, n702_o, n699_o, n696_o, n693_o, n690_o, n687_o, n684_o, n681_o, n678_o, n675_o, n672_o, n669_o, n666_o, n663_o, n660_o, n657_o, n654_o, n651_o, n648_o, n645_o, n642_o, n639_o, n636_o, n633_o, n630_o, n627_o, n624_o, n621_o, n618_o, n615_o, n612_o, n609_o, n606_o, n603_o, n600_o, n597_o, n594_o, n591_o, n588_o, n585_o, n582_o, n579_o, n576_o, n573_o, n570_o, n567_o, n564_o, n561_o, n558_o, n555_o, n552_o, n549_o, n546_o, n543_o, n540_o, n537_o, n534_o, n531_o, n528_o, n525_o, n522_o, n519_o, n516_o, n513_o, n510_o, n507_o, n504_o, n501_o, n498_o, n495_o, n492_o, n489_o, n486_o, n483_o, n480_o, n477_o, n474_o, n471_o, n468_o, n465_o, n462_o, n459_o, n456_o, n453_o, n450_o, n447_o, n444_o, n441_o, n438_o, n435_o, n432_o, n429_o, n426_o, n423_o, n420_o, n417_o, n414_o, n411_o, n408_o, n405_o, n402_o, n399_o, n396_o, n393_o, n390_o, n387_o, n384_o, n381_o, n378_o, n375_o, n372_o, n369_o, n366_o, n363_o, n360_o, n357_o, n354_o, n351_o, n348_o, n345_o, n342_o, n339_o, n336_o, n333_o, n330_o, n327_o, n324_o, n321_o, n318_o, n315_o, n312_o, n309_o, n306_o, n303_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:35:4  */
    always @*
        case (n1838_o)
            512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n1839_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n1839_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n1839_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n1839_o = 3'b000;
            default: n1839_o = 3'bXXX;
        endcase
endmodule

module fdiv#(parameter ID=1)
    (input wire clk,
        input wire[10:0] X,
        input wire[10:0] Y,
        output wire[10:0] R);
    wire[4:0] fx;
    wire[4:0] fy;
    wire[5:0] expr0;
    wire[5:0] expr0_d1;
    wire[5:0] expr0_d2;
    wire[5:0] expr0_d3;
    wire sr;
    wire sr_d1;
    wire sr_d2;
    wire sr_d3;
    wire[3:0] exnxy;
    wire[1:0] exnr0;
    wire[1:0] exnr0_d1;
    wire[1:0] exnr0_d2;
    wire[1:0] exnr0_d3;
    wire[4:0] d;
    wire[4:0] d_d1;
    wire[4:0] d_d2;
    wire[5:0] psx;
    wire[7:0] betaw4;
    wire[8:0] sel4;
    wire[2:0] q4;
    wire[2:0] q4_copy5;
    wire[7:0] absq4d;
    wire[7:0] w3;
    wire[7:0] betaw3;
    wire[7:0] betaw3_d1;
    wire[8:0] sel3;
    wire[2:0] q3;
    wire[2:0] q3_copy6;
    wire[2:0] q3_copy6_d1;
    wire[7:0] absq3d;
    wire[7:0] w2;
    wire[7:0] betaw2;
    wire[7:0] betaw2_d1;
    wire[8:0] sel2;
    wire[2:0] q2;
    wire[2:0] q2_copy7;
    wire[2:0] q2_copy7_d1;
    wire[7:0] absq2d;
    wire[7:0] w1;
    wire[7:0] betaw1;
    wire[7:0] betaw1_d1;
    wire[8:0] sel1;
    wire[2:0] q1;
    wire[2:0] q1_d1;
    wire[2:0] q1_copy8;
    wire[7:0] absq1d;
    wire[7:0] absq1d_d1;
    wire[7:0] w0;
    wire[5:0] wfinal;
    wire qm0;
    wire[1:0] qp4;
    wire[1:0] qp4_d1;
    wire[1:0] qp4_d2;
    wire[1:0] qm4;
    wire[1:0] qm4_d1;
    wire[1:0] qm4_d2;
    wire[1:0] qm4_d3;
    wire[1:0] qp3;
    wire[1:0] qp3_d1;
    wire[1:0] qm3;
    wire[1:0] qm3_d1;
    wire[1:0] qm3_d2;
    wire[1:0] qp2;
    wire[1:0] qm2;
    wire[1:0] qm2_d1;
    wire[1:0] qp1;
    wire[1:0] qm1;
    wire[1:0] qm1_d1;
    wire[7:0] qp;
    wire[7:0] qp_d1;
    wire[7:0] qm;
    wire[7:0] quotient;
    wire[6:0] mr;
    wire[4:0] frnorm;
    wire round;
    wire[5:0] expr1;
    wire[9:0] expfrac;
    wire[9:0] expfracr;
    wire[1:0] exnr;
    wire[1:0] exnrfinal;
    wire[3:0] n34_o;
    wire[4:0] n36_o;
    wire[3:0] n37_o;
    wire[4:0] n39_o;
    wire[3:0] n40_o;
    wire[5:0] n42_o;
    wire[3:0] n43_o;
    wire[5:0] n45_o;
    wire[5:0] n46_o;
    wire n47_o;
    wire n48_o;
    wire n49_o;
    wire[1:0] n50_o;
    wire[1:0] n51_o;
    wire[3:0] n52_o;
    wire n55_o;
    wire n58_o;
    wire n60_o;
    wire n61_o;
    wire n63_o;
    wire n64_o;
    wire n67_o;
    wire n69_o;
    wire n70_o;
    wire n72_o;
    wire n73_o;
    wire[2:0] n75_o;
    reg[1:0] n76_o;
    wire[5:0] n78_o;
    wire[7:0] n80_o;
    wire[5:0] n81_o;
    wire[2:0] n82_o;
    wire[8:0] n83_o;
    wire[2:0] selfunctiontable4_n84;
    wire[2:0] selfunctiontable4_y;
    wire[7:0] n88_o;
    wire n90_o;
    wire n92_o;
    wire n93_o;
    wire[6:0] n95_o;
    wire[7:0] n97_o;
    wire n99_o;
    wire n101_o;
    wire n102_o;
    wire[1:0] n104_o;
    reg[7:0] n105_o;
    wire n106_o;
    wire[7:0] n107_o;
    wire n109_o;
    wire[7:0] n110_o;
    reg[7:0] n111_o;
    wire[5:0] n112_o;
    wire[7:0] n114_o;
    wire[5:0] n115_o;
    wire[2:0] n116_o;
    wire[8:0] n117_o;
    wire[2:0] selfunctiontable3_n118;
    wire[2:0] selfunctiontable3_y;
    wire[7:0] n122_o;
    wire n124_o;
    wire n126_o;
    wire n127_o;
    wire[6:0] n129_o;
    wire[7:0] n131_o;
    wire n133_o;
    wire n135_o;
    wire n136_o;
    wire[1:0] n138_o;
    reg[7:0] n139_o;
    wire n140_o;
    wire[7:0] n141_o;
    wire n143_o;
    wire[7:0] n144_o;
    reg[7:0] n145_o;
    wire[5:0] n146_o;
    wire[7:0] n148_o;
    wire[5:0] n149_o;
    wire[2:0] n150_o;
    wire[8:0] n151_o;
    wire[2:0] selfunctiontable2_n152;
    wire[2:0] selfunctiontable2_y;
    wire[7:0] n156_o;
    wire n158_o;
    wire n160_o;
    wire n161_o;
    wire[6:0] n163_o;
    wire[7:0] n165_o;
    wire n167_o;
    wire n169_o;
    wire n170_o;
    wire[1:0] n172_o;
    reg[7:0] n173_o;
    wire n174_o;
    wire[7:0] n175_o;
    wire n177_o;
    wire[7:0] n178_o;
    reg[7:0] n179_o;
    wire[5:0] n180_o;
    wire[7:0] n182_o;
    wire[5:0] n183_o;
    wire[2:0] n184_o;
    wire[8:0] n185_o;
    wire[2:0] selfunctiontable1_n186;
    wire[2:0] selfunctiontable1_y;
    wire[7:0] n190_o;
    wire n192_o;
    wire n194_o;
    wire n195_o;
    wire[6:0] n197_o;
    wire[7:0] n199_o;
    wire n201_o;
    wire n203_o;
    wire n204_o;
    wire[1:0] n206_o;
    reg[7:0] n207_o;
    wire n208_o;
    wire[7:0] n209_o;
    wire n211_o;
    wire[7:0] n212_o;
    reg[7:0] n213_o;
    wire[5:0] n214_o;
    wire n215_o;
    wire[1:0] n216_o;
    wire n217_o;
    wire[1:0] n219_o;
    wire[1:0] n220_o;
    wire n221_o;
    wire[1:0] n223_o;
    wire[1:0] n224_o;
    wire n225_o;
    wire[1:0] n227_o;
    wire[1:0] n228_o;
    wire n229_o;
    wire[1:0] n231_o;
    wire[3:0] n232_o;
    wire[5:0] n233_o;
    wire[7:0] n234_o;
    wire n235_o;
    wire[2:0] n236_o;
    wire[4:0] n237_o;
    wire[6:0] n238_o;
    wire[7:0] n239_o;
    wire[7:0] n240_o;
    wire[6:0] n241_o;
    wire[4:0] n242_o;
    wire n243_o;
    wire[4:0] n244_o;
    wire[4:0] n245_o;
    wire n246_o;
    wire n247_o;
    wire[5:0] n249_o;
    wire[5:0] n250_o;
    wire[3:0] n251_o;
    wire[9:0] n252_o;
    wire[9:0] n254_o;
    wire[9:0] n255_o;
    wire n257_o;
    wire[1:0] n258_o;
    wire[1:0] n260_o;
    wire n262_o;
    wire[1:0] n263_o;
    wire n266_o;
    reg[1:0] n267_o;
    wire[2:0] n268_o;
    wire[7:0] n269_o;
    wire[10:0] n270_o;
    reg[5:0] n271_q;
    reg[5:0] n272_q;
    reg[5:0] n273_q;
    reg n274_q;
    reg n275_q;
    reg n276_q;
    reg[1:0] n277_q;
    reg[1:0] n278_q;
    reg[1:0] n279_q;
    reg[4:0] n280_q;
    reg[4:0] n281_q;
    reg[7:0] n282_q;
    reg[2:0] n283_q;
    reg[7:0] n284_q;
    reg[2:0] n285_q;
    reg[7:0] n286_q;
    reg[2:0] n287_q;
    reg[7:0] n288_q;
    reg[1:0] n289_q;
    reg[1:0] n290_q;
    reg[1:0] n291_q;
    reg[1:0] n292_q;
    reg[1:0] n293_q;
    reg[1:0] n294_q;
    reg[1:0] n295_q;
    reg[1:0] n296_q;
    reg[1:0] n297_q;
    reg[1:0] n298_q;
    reg[7:0] n299_q;
    assign R = n270_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:588:8  */
    assign fx = n36_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:589:8  */
    assign fy = n39_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:590:8  */
    assign expr0 = n46_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:590:15  */
    assign expr0_d1 = n271_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:590:25  */
    assign expr0_d2 = n272_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:590:35  */
    assign expr0_d3 = n273_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:591:8  */
    assign sr = n49_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:591:12  */
    assign sr_d1 = n274_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:591:19  */
    assign sr_d2 = n275_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:591:26  */
    assign sr_d3 = n276_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:592:8  */
    assign exnxy = n52_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:593:8  */
    assign exnr0 = n76_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:593:15  */
    assign exnr0_d1 = n277_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:593:25  */
    assign exnr0_d2 = n278_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:593:35  */
    assign exnr0_d3 = n279_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:594:8  */
    assign d = fy; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:594:11  */
    assign d_d1 = n280_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:594:17  */
    assign d_d2 = n281_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:595:8  */
    assign psx = n78_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:596:8  */
    assign betaw4 = n80_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:597:8  */
    assign sel4 = n83_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:598:8  */
    assign q4 = q4_copy5; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:599:8  */
    assign q4_copy5 = selfunctiontable4_n84; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:600:8  */
    assign absq4d = n105_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:601:8  */
    assign w3 = n111_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:602:8  */
    assign betaw3 = n114_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:602:16  */
    assign betaw3_d1 = n282_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:603:8  */
    assign sel3 = n117_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:604:8  */
    assign q3 = q3_copy6_d1; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:605:8  */
    assign q3_copy6 = selfunctiontable3_n118; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:605:18  */
    assign q3_copy6_d1 = n283_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:606:8  */
    assign absq3d = n139_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:607:8  */
    assign w2 = n145_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:608:8  */
    assign betaw2 = n148_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:608:16  */
    assign betaw2_d1 = n284_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:609:8  */
    assign sel2 = n151_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:610:8  */
    assign q2 = q2_copy7_d1; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:611:8  */
    assign q2_copy7 = selfunctiontable2_n152; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:611:18  */
    assign q2_copy7_d1 = n285_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:612:8  */
    assign absq2d = n173_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:613:8  */
    assign w1 = n179_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:614:8  */
    assign betaw1 = n182_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:614:16  */
    assign betaw1_d1 = n286_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:615:8  */
    assign sel1 = n185_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:616:8  */
    assign q1 = q1_copy8; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:616:12  */
    assign q1_d1 = n287_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:617:8  */
    assign q1_copy8 = selfunctiontable1_n186; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:618:8  */
    assign absq1d = n207_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:618:16  */
    assign absq1d_d1 = n288_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:619:8  */
    assign w0 = n213_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:620:8  */
    assign wfinal = n214_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:621:8  */
    assign qm0 = n215_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:622:8  */
    assign qp4 = n216_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:622:13  */
    assign qp4_d1 = n289_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:622:21  */
    assign qp4_d2 = n290_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:623:8  */
    assign qm4 = n219_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:623:13  */
    assign qm4_d1 = n291_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:623:21  */
    assign qm4_d2 = n292_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:623:29  */
    assign qm4_d3 = n293_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:624:8  */
    assign qp3 = n220_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:624:13  */
    assign qp3_d1 = n294_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:625:8  */
    assign qm3 = n223_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:625:13  */
    assign qm3_d1 = n295_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:625:21  */
    assign qm3_d2 = n296_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:626:8  */
    assign qp2 = n224_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:627:8  */
    assign qm2 = n227_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:627:13  */
    assign qm2_d1 = n297_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:628:8  */
    assign qp1 = n228_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:629:8  */
    assign qm1 = n231_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:629:13  */
    assign qm1_d1 = n298_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:630:8  */
    assign qp = n234_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:630:12  */
    assign qp_d1 = n299_q; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:631:8  */
    assign qm = n239_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:632:8  */
    assign quotient = n240_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:633:8  */
    assign mr = n241_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:634:8  */
    assign frnorm = n244_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:635:8  */
    assign round = n246_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:636:8  */
    assign expr1 = n250_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:637:8  */
    assign expfrac = n252_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:638:8  */
    assign expfracr = n255_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:639:8  */
    assign exnr = n258_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:640:8  */
    assign exnrfinal = n267_o; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:676:17  */
    assign n34_o = X[3:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:676:14  */
    assign n36_o = {1'b1, n34_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:677:17  */
    assign n37_o = Y[3:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:677:14  */
    assign n39_o = {1'b1, n37_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:679:22  */
    assign n40_o = X[7:4];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:679:19  */
    assign n42_o = {2'b00, n40_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:679:47  */
    assign n43_o = Y[7:4];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:679:44  */
    assign n45_o = {2'b00, n43_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:679:36  */
    assign n46_o = n42_o-n45_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:680:11  */
    assign n47_o = X[8];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:680:20  */
    assign n48_o = Y[8];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:680:15  */
    assign n49_o = n47_o ^ n48_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:682:14  */
    assign n50_o = X[10:9];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:682:31  */
    assign n51_o = Y[10:9];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:682:28  */
    assign n52_o = {n50_o, n51_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:685:18  */
    assign n55_o = exnxy == 4'b0101;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:686:18  */
    assign n58_o = exnxy == 4'b0001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:686:30  */
    assign n60_o = exnxy == 4'b0010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:686:30  */
    assign n61_o = n58_o | n60_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:686:39  */
    assign n63_o = exnxy == 4'b0110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:686:39  */
    assign n64_o = n61_o | n63_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:687:18  */
    assign n67_o = exnxy == 4'b0100;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:687:30  */
    assign n69_o = exnxy == 4'b1000;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:687:30  */
    assign n70_o = n67_o | n69_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:687:39  */
    assign n72_o = exnxy == 4'b1001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:687:39  */
    assign n73_o = n70_o | n72_o;
    assign n75_o = {n73_o, n64_o, n55_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:683:4  */
    always @*
        case (n75_o)
            3'b100: n76_o = 2'b10;
            3'b010: n76_o = 2'b00;
            3'b001: n76_o = 2'b01;
            default: n76_o = 2'b11;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:690:15  */
    assign n78_o = {1'b0, fx};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:691:20  */
    assign n80_o = {2'b00, psx};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:692:18  */
    assign n81_o = betaw4[7:2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:692:34  */
    assign n82_o = d[3:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:692:31  */
    assign n83_o = {n81_o, n82_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:695:23  */
    assign selfunctiontable4_n84 = selfunctiontable4_y; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:693:4  */
    selfunction_f300_uid4 selfunctiontable4(
        .x(sel4),
        .y(selfunctiontable4_y));
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:700:16  */
    assign n88_o = {3'b000, d};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:700:66  */
    assign n90_o = q4 == 3'b001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:700:77  */
    assign n92_o = q4 == 3'b111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:700:77  */
    assign n93_o = n90_o | n92_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:701:15  */
    assign n95_o = {2'b00, d};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:701:19  */
    assign n97_o = {n95_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:701:52  */
    assign n99_o = q4 == 3'b010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:701:63  */
    assign n101_o = q4 == 3'b110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:701:63  */
    assign n102_o = n99_o | n101_o;
    assign n104_o = {n102_o, n93_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:698:4  */
    always @*
        case (n104_o)
            2'b10: n105_o = n97_o;
            2'b01: n105_o = n88_o;
            default: n105_o = 8'b00000000;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:704:11  */
    assign n106_o = q4[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:705:16  */
    assign n107_o = betaw4-absq4d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:705:25  */
    assign n109_o = n106_o == 1'b0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:706:17  */
    assign n110_o = betaw4+absq4d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:704:4  */
    always @*
        case (n109_o)
            1'b1: n111_o = n107_o;
            default: n111_o = n110_o;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:708:16  */
    assign n112_o = w3[5:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:708:29  */
    assign n114_o = {n112_o, 2'b00};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:709:18  */
    assign n115_o = betaw3[7:2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:709:34  */
    assign n116_o = d[3:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:709:31  */
    assign n117_o = {n115_o, n116_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:712:23  */
    assign selfunctiontable3_n118 = selfunctiontable3_y; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:710:4  */
    selfunction_f300_uid4 selfunctiontable3(
        .x(sel3),
        .y(selfunctiontable3_y));
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:717:16  */
    assign n122_o = {3'b000, d_d1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:717:66  */
    assign n124_o = q3 == 3'b001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:717:77  */
    assign n126_o = q3 == 3'b111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:717:77  */
    assign n127_o = n124_o | n126_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:718:15  */
    assign n129_o = {2'b00, d_d1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:718:22  */
    assign n131_o = {n129_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:718:52  */
    assign n133_o = q3 == 3'b010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:718:63  */
    assign n135_o = q3 == 3'b110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:718:63  */
    assign n136_o = n133_o | n135_o;
    assign n138_o = {n136_o, n127_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:715:4  */
    always @*
        case (n138_o)
            2'b10: n139_o = n131_o;
            2'b01: n139_o = n122_o;
            default: n139_o = 8'b00000000;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:721:11  */
    assign n140_o = q3[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:722:19  */
    assign n141_o = betaw3_d1-absq3d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:722:28  */
    assign n143_o = n140_o == 1'b0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:723:20  */
    assign n144_o = betaw3_d1+absq3d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:721:4  */
    always @*
        case (n143_o)
            1'b1: n145_o = n141_o;
            default: n145_o = n144_o;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:725:16  */
    assign n146_o = w2[5:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:725:29  */
    assign n148_o = {n146_o, 2'b00};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:726:18  */
    assign n149_o = betaw2[7:2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:726:37  */
    assign n150_o = d_d1[3:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:726:31  */
    assign n151_o = {n149_o, n150_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:729:23  */
    assign selfunctiontable2_n152 = selfunctiontable2_y; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:727:4  */
    selfunction_f300_uid4 selfunctiontable2(
        .x(sel2),
        .y(selfunctiontable2_y));
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:734:16  */
    assign n156_o = {3'b000, d_d2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:734:66  */
    assign n158_o = q2 == 3'b001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:734:77  */
    assign n160_o = q2 == 3'b111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:734:77  */
    assign n161_o = n158_o | n160_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:735:15  */
    assign n163_o = {2'b00, d_d2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:735:22  */
    assign n165_o = {n163_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:735:52  */
    assign n167_o = q2 == 3'b010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:735:63  */
    assign n169_o = q2 == 3'b110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:735:63  */
    assign n170_o = n167_o | n169_o;
    assign n172_o = {n170_o, n161_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:732:4  */
    always @*
        case (n172_o)
            2'b10: n173_o = n165_o;
            2'b01: n173_o = n156_o;
            default: n173_o = 8'b00000000;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:738:11  */
    assign n174_o = q2[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:739:19  */
    assign n175_o = betaw2_d1-absq2d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:739:28  */
    assign n177_o = n174_o == 1'b0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:740:20  */
    assign n178_o = betaw2_d1+absq2d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:738:4  */
    always @*
        case (n177_o)
            1'b1: n179_o = n175_o;
            default: n179_o = n178_o;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:742:16  */
    assign n180_o = w1[5:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:742:29  */
    assign n182_o = {n180_o, 2'b00};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:743:18  */
    assign n183_o = betaw1[7:2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:743:37  */
    assign n184_o = d_d2[3:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:743:31  */
    assign n185_o = {n183_o, n184_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:746:23  */
    assign selfunctiontable1_n186 = selfunctiontable1_y; // (signal)
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:744:4  */
    selfunction_f300_uid4 selfunctiontable1(
        .x(sel1),
        .y(selfunctiontable1_y));
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:751:16  */
    assign n190_o = {3'b000, d_d2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:751:66  */
    assign n192_o = q1 == 3'b001;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:751:77  */
    assign n194_o = q1 == 3'b111;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:751:77  */
    assign n195_o = n192_o | n194_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:752:15  */
    assign n197_o = {2'b00, d_d2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:752:22  */
    assign n199_o = {n197_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:752:52  */
    assign n201_o = q1 == 3'b010;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:752:63  */
    assign n203_o = q1 == 3'b110;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:752:63  */
    assign n204_o = n201_o | n203_o;
    assign n206_o = {n204_o, n195_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:749:4  */
    always @*
        case (n206_o)
            2'b10: n207_o = n199_o;
            2'b01: n207_o = n190_o;
            default: n207_o = 8'b00000000;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:755:14  */
    assign n208_o = q1_d1[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:756:19  */
    assign n209_o = betaw1_d1-absq1d_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:756:31  */
    assign n211_o = n208_o == 1'b0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:757:20  */
    assign n212_o = betaw1_d1+absq1d_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:755:4  */
    always @*
        case (n211_o)
            1'b1: n213_o = n209_o;
            default: n213_o = n212_o;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:759:16  */
    assign n214_o = w0[5:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:760:17  */
    assign n215_o = wfinal[5];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:761:18  */
    assign n216_o = q4[1:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:762:18  */
    assign n217_o = q4[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:762:22  */
    assign n219_o = {n217_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:763:18  */
    assign n220_o = q3[1:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:764:18  */
    assign n221_o = q3[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:764:22  */
    assign n223_o = {n221_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:765:18  */
    assign n224_o = q2[1:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:766:18  */
    assign n225_o = q2[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:766:22  */
    assign n227_o = {n225_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:767:18  */
    assign n228_o = q1[1:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:768:18  */
    assign n229_o = q1[2];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:768:22  */
    assign n231_o = {n229_o, 1'b0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:769:17  */
    assign n232_o = {qp4_d2, qp3_d1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:769:26  */
    assign n233_o = {n232_o, qp2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:769:32  */
    assign n234_o = {n233_o, qp1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:770:16  */
    assign n235_o = qm4_d3[0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:770:20  */
    assign n236_o = {n235_o, qm3_d2};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:770:29  */
    assign n237_o = {n236_o, qm2_d1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:770:38  */
    assign n238_o = {n237_o, qm1_d1};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:770:47  */
    assign n239_o = {n238_o, qm0};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:771:22  */
    assign n240_o = qp_d1-qm;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:775:18  */
    assign n241_o = quotient[6:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:777:19  */
    assign n242_o = mr[5:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:777:40  */
    assign n243_o = mr[6];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:777:33  */
    assign n244_o = n243_o ? n242_o : n245_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:778:19  */
    assign n245_o = mr[4:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:779:19  */
    assign n246_o = frnorm[0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:780:57  */
    assign n247_o = mr[6];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:780:53  */
    assign n249_o = {5'b00011, n247_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:780:22  */
    assign n250_o = expr0_d3+n249_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:782:29  */
    assign n251_o = frnorm[4:1];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:782:21  */
    assign n252_o = {expr1, n251_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:783:47  */
    assign n254_o = {9'b000000000, round};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:783:24  */
    assign n255_o = expfrac+n254_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:784:36  */
    assign n257_o = expfracr[9];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:784:23  */
    assign n258_o = n257_o ? 2'b00 : n263_o;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:785:37  */
    assign n260_o = expfracr[9:8];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:785:50  */
    assign n262_o = n260_o == 2'b01;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:785:12  */
    assign n263_o = n262_o ? 2'b10 : 2'b01;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:789:17  */
    assign n266_o = exnr0_d3 == 2'b01;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:787:4  */
    always @*
        case (n266_o)
            1'b1: n267_o = exnr;
            default: n267_o = exnr0_d3;
        endcase
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:791:19  */
    assign n268_o = {exnrfinal, sr_d3};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:791:37  */
    assign n269_o = expfracr[7:0];
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:791:27  */
    assign n270_o = {n268_o, n269_o};
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n271_q <= expr0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n272_q <= expr0_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n273_q <= expr0_d2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n274_q <= sr;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n275_q <= sr_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n276_q <= sr_d2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n277_q <= exnr0;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n278_q <= exnr0_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n279_q <= exnr0_d2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n280_q <= d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n281_q <= d_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n282_q <= betaw3;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n283_q <= q3_copy6;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n284_q <= betaw2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n285_q <= q2_copy7;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n286_q <= betaw1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n287_q <= q1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n288_q <= absq1d;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n289_q <= qp4;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n290_q <= qp4_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n291_q <= qm4;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n292_q <= qm4_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n293_q <= qm4_d2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n294_q <= qp3;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n295_q <= qm3;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n296_q <= qm3_d1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n297_q <= qm2;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n298_q <= qm1;
    /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_4.vhdl:644:10  */
    always @(posedge clk)
        n299_q <= qp;
endmodule

