module selfunction_f300_uid4
  (input  [8:0] x,
   output [2:0] y);
  wire [2:0] y0;
  wire [2:0] y1;
  wire n1127_o;
  wire n1130_o;
  wire n1133_o;
  wire n1136_o;
  wire n1139_o;
  wire n1142_o;
  wire n1145_o;
  wire n1148_o;
  wire n1151_o;
  wire n1154_o;
  wire n1157_o;
  wire n1160_o;
  wire n1163_o;
  wire n1166_o;
  wire n1169_o;
  wire n1172_o;
  wire n1175_o;
  wire n1178_o;
  wire n1181_o;
  wire n1184_o;
  wire n1187_o;
  wire n1190_o;
  wire n1193_o;
  wire n1196_o;
  wire n1199_o;
  wire n1202_o;
  wire n1205_o;
  wire n1208_o;
  wire n1211_o;
  wire n1214_o;
  wire n1217_o;
  wire n1220_o;
  wire n1223_o;
  wire n1226_o;
  wire n1229_o;
  wire n1232_o;
  wire n1235_o;
  wire n1238_o;
  wire n1241_o;
  wire n1244_o;
  wire n1247_o;
  wire n1250_o;
  wire n1253_o;
  wire n1256_o;
  wire n1259_o;
  wire n1262_o;
  wire n1265_o;
  wire n1268_o;
  wire n1271_o;
  wire n1274_o;
  wire n1277_o;
  wire n1280_o;
  wire n1283_o;
  wire n1286_o;
  wire n1289_o;
  wire n1292_o;
  wire n1295_o;
  wire n1298_o;
  wire n1301_o;
  wire n1304_o;
  wire n1307_o;
  wire n1310_o;
  wire n1313_o;
  wire n1316_o;
  wire n1319_o;
  wire n1322_o;
  wire n1325_o;
  wire n1328_o;
  wire n1331_o;
  wire n1334_o;
  wire n1337_o;
  wire n1340_o;
  wire n1343_o;
  wire n1346_o;
  wire n1349_o;
  wire n1352_o;
  wire n1355_o;
  wire n1358_o;
  wire n1361_o;
  wire n1364_o;
  wire n1367_o;
  wire n1370_o;
  wire n1373_o;
  wire n1376_o;
  wire n1379_o;
  wire n1382_o;
  wire n1385_o;
  wire n1388_o;
  wire n1391_o;
  wire n1394_o;
  wire n1397_o;
  wire n1400_o;
  wire n1403_o;
  wire n1406_o;
  wire n1409_o;
  wire n1412_o;
  wire n1415_o;
  wire n1418_o;
  wire n1421_o;
  wire n1424_o;
  wire n1427_o;
  wire n1430_o;
  wire n1433_o;
  wire n1436_o;
  wire n1439_o;
  wire n1442_o;
  wire n1445_o;
  wire n1448_o;
  wire n1451_o;
  wire n1454_o;
  wire n1457_o;
  wire n1460_o;
  wire n1463_o;
  wire n1466_o;
  wire n1469_o;
  wire n1472_o;
  wire n1475_o;
  wire n1478_o;
  wire n1481_o;
  wire n1484_o;
  wire n1487_o;
  wire n1490_o;
  wire n1493_o;
  wire n1496_o;
  wire n1499_o;
  wire n1502_o;
  wire n1505_o;
  wire n1508_o;
  wire n1511_o;
  wire n1514_o;
  wire n1517_o;
  wire n1520_o;
  wire n1523_o;
  wire n1526_o;
  wire n1529_o;
  wire n1532_o;
  wire n1535_o;
  wire n1538_o;
  wire n1541_o;
  wire n1544_o;
  wire n1547_o;
  wire n1550_o;
  wire n1553_o;
  wire n1556_o;
  wire n1559_o;
  wire n1562_o;
  wire n1565_o;
  wire n1568_o;
  wire n1571_o;
  wire n1574_o;
  wire n1577_o;
  wire n1580_o;
  wire n1583_o;
  wire n1586_o;
  wire n1589_o;
  wire n1592_o;
  wire n1595_o;
  wire n1598_o;
  wire n1601_o;
  wire n1604_o;
  wire n1607_o;
  wire n1610_o;
  wire n1613_o;
  wire n1616_o;
  wire n1619_o;
  wire n1622_o;
  wire n1625_o;
  wire n1628_o;
  wire n1631_o;
  wire n1634_o;
  wire n1637_o;
  wire n1640_o;
  wire n1643_o;
  wire n1646_o;
  wire n1649_o;
  wire n1652_o;
  wire n1655_o;
  wire n1658_o;
  wire n1661_o;
  wire n1664_o;
  wire n1667_o;
  wire n1670_o;
  wire n1673_o;
  wire n1676_o;
  wire n1679_o;
  wire n1682_o;
  wire n1685_o;
  wire n1688_o;
  wire n1691_o;
  wire n1694_o;
  wire n1697_o;
  wire n1700_o;
  wire n1703_o;
  wire n1706_o;
  wire n1709_o;
  wire n1712_o;
  wire n1715_o;
  wire n1718_o;
  wire n1721_o;
  wire n1724_o;
  wire n1727_o;
  wire n1730_o;
  wire n1733_o;
  wire n1736_o;
  wire n1739_o;
  wire n1742_o;
  wire n1745_o;
  wire n1748_o;
  wire n1751_o;
  wire n1754_o;
  wire n1757_o;
  wire n1760_o;
  wire n1763_o;
  wire n1766_o;
  wire n1769_o;
  wire n1772_o;
  wire n1775_o;
  wire n1778_o;
  wire n1781_o;
  wire n1784_o;
  wire n1787_o;
  wire n1790_o;
  wire n1793_o;
  wire n1796_o;
  wire n1799_o;
  wire n1802_o;
  wire n1805_o;
  wire n1808_o;
  wire n1811_o;
  wire n1814_o;
  wire n1817_o;
  wire n1820_o;
  wire n1823_o;
  wire n1826_o;
  wire n1829_o;
  wire n1832_o;
  wire n1835_o;
  wire n1838_o;
  wire n1841_o;
  wire n1844_o;
  wire n1847_o;
  wire n1850_o;
  wire n1853_o;
  wire n1856_o;
  wire n1859_o;
  wire n1862_o;
  wire n1865_o;
  wire n1868_o;
  wire n1871_o;
  wire n1874_o;
  wire n1877_o;
  wire n1880_o;
  wire n1883_o;
  wire n1886_o;
  wire n1889_o;
  wire n1892_o;
  wire n1895_o;
  wire n1898_o;
  wire n1901_o;
  wire n1904_o;
  wire n1907_o;
  wire n1910_o;
  wire n1913_o;
  wire n1916_o;
  wire n1919_o;
  wire n1922_o;
  wire n1925_o;
  wire n1928_o;
  wire n1931_o;
  wire n1934_o;
  wire n1937_o;
  wire n1940_o;
  wire n1943_o;
  wire n1946_o;
  wire n1949_o;
  wire n1952_o;
  wire n1955_o;
  wire n1958_o;
  wire n1961_o;
  wire n1964_o;
  wire n1967_o;
  wire n1970_o;
  wire n1973_o;
  wire n1976_o;
  wire n1979_o;
  wire n1982_o;
  wire n1985_o;
  wire n1988_o;
  wire n1991_o;
  wire n1994_o;
  wire n1997_o;
  wire n2000_o;
  wire n2003_o;
  wire n2006_o;
  wire n2009_o;
  wire n2012_o;
  wire n2015_o;
  wire n2018_o;
  wire n2021_o;
  wire n2024_o;
  wire n2027_o;
  wire n2030_o;
  wire n2033_o;
  wire n2036_o;
  wire n2039_o;
  wire n2042_o;
  wire n2045_o;
  wire n2048_o;
  wire n2051_o;
  wire n2054_o;
  wire n2057_o;
  wire n2060_o;
  wire n2063_o;
  wire n2066_o;
  wire n2069_o;
  wire n2072_o;
  wire n2075_o;
  wire n2078_o;
  wire n2081_o;
  wire n2084_o;
  wire n2087_o;
  wire n2090_o;
  wire n2093_o;
  wire n2096_o;
  wire n2099_o;
  wire n2102_o;
  wire n2105_o;
  wire n2108_o;
  wire n2111_o;
  wire n2114_o;
  wire n2117_o;
  wire n2120_o;
  wire n2123_o;
  wire n2126_o;
  wire n2129_o;
  wire n2132_o;
  wire n2135_o;
  wire n2138_o;
  wire n2141_o;
  wire n2144_o;
  wire n2147_o;
  wire n2150_o;
  wire n2153_o;
  wire n2156_o;
  wire n2159_o;
  wire n2162_o;
  wire n2165_o;
  wire n2168_o;
  wire n2171_o;
  wire n2174_o;
  wire n2177_o;
  wire n2180_o;
  wire n2183_o;
  wire n2186_o;
  wire n2189_o;
  wire n2192_o;
  wire n2195_o;
  wire n2198_o;
  wire n2201_o;
  wire n2204_o;
  wire n2207_o;
  wire n2210_o;
  wire n2213_o;
  wire n2216_o;
  wire n2219_o;
  wire n2222_o;
  wire n2225_o;
  wire n2228_o;
  wire n2231_o;
  wire n2234_o;
  wire n2237_o;
  wire n2240_o;
  wire n2243_o;
  wire n2246_o;
  wire n2249_o;
  wire n2252_o;
  wire n2255_o;
  wire n2258_o;
  wire n2261_o;
  wire n2264_o;
  wire n2267_o;
  wire n2270_o;
  wire n2273_o;
  wire n2276_o;
  wire n2279_o;
  wire n2282_o;
  wire n2285_o;
  wire n2288_o;
  wire n2291_o;
  wire n2294_o;
  wire n2297_o;
  wire n2300_o;
  wire n2303_o;
  wire n2306_o;
  wire n2309_o;
  wire n2312_o;
  wire n2315_o;
  wire n2318_o;
  wire n2321_o;
  wire n2324_o;
  wire n2327_o;
  wire n2330_o;
  wire n2333_o;
  wire n2336_o;
  wire n2339_o;
  wire n2342_o;
  wire n2345_o;
  wire n2348_o;
  wire n2351_o;
  wire n2354_o;
  wire n2357_o;
  wire n2360_o;
  wire n2363_o;
  wire n2366_o;
  wire n2369_o;
  wire n2372_o;
  wire n2375_o;
  wire n2378_o;
  wire n2381_o;
  wire n2384_o;
  wire n2387_o;
  wire n2390_o;
  wire n2393_o;
  wire n2396_o;
  wire n2399_o;
  wire n2402_o;
  wire n2405_o;
  wire n2408_o;
  wire n2411_o;
  wire n2414_o;
  wire n2417_o;
  wire n2420_o;
  wire n2423_o;
  wire n2426_o;
  wire n2429_o;
  wire n2432_o;
  wire n2435_o;
  wire n2438_o;
  wire n2441_o;
  wire n2444_o;
  wire n2447_o;
  wire n2450_o;
  wire n2453_o;
  wire n2456_o;
  wire n2459_o;
  wire n2462_o;
  wire n2465_o;
  wire n2468_o;
  wire n2471_o;
  wire n2474_o;
  wire n2477_o;
  wire n2480_o;
  wire n2483_o;
  wire n2486_o;
  wire n2489_o;
  wire n2492_o;
  wire n2495_o;
  wire n2498_o;
  wire n2501_o;
  wire n2504_o;
  wire n2507_o;
  wire n2510_o;
  wire n2513_o;
  wire n2516_o;
  wire n2519_o;
  wire n2522_o;
  wire n2525_o;
  wire n2528_o;
  wire n2531_o;
  wire n2534_o;
  wire n2537_o;
  wire n2540_o;
  wire n2543_o;
  wire n2546_o;
  wire n2549_o;
  wire n2552_o;
  wire n2555_o;
  wire n2558_o;
  wire n2561_o;
  wire n2564_o;
  wire n2567_o;
  wire n2570_o;
  wire n2573_o;
  wire n2576_o;
  wire n2579_o;
  wire n2582_o;
  wire n2585_o;
  wire n2588_o;
  wire n2591_o;
  wire n2594_o;
  wire n2597_o;
  wire n2600_o;
  wire n2603_o;
  wire n2606_o;
  wire n2609_o;
  wire n2612_o;
  wire n2615_o;
  wire n2618_o;
  wire n2621_o;
  wire n2624_o;
  wire n2627_o;
  wire n2630_o;
  wire n2633_o;
  wire n2636_o;
  wire n2639_o;
  wire n2642_o;
  wire n2645_o;
  wire n2648_o;
  wire n2651_o;
  wire n2654_o;
  wire n2657_o;
  wire n2660_o;
  wire [511:0] n2662_o;
  reg [2:0] n2663_o;
  assign y = y1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:28:8  */
  assign y0 = n2663_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:33:8  */
  assign y1 = y0; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:36:13  */
  assign n1127_o = x == 9'b000000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:37:13  */
  assign n1130_o = x == 9'b000000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:38:13  */
  assign n1133_o = x == 9'b000000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:39:13  */
  assign n1136_o = x == 9'b000000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:40:13  */
  assign n1139_o = x == 9'b000000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:41:13  */
  assign n1142_o = x == 9'b000000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:42:13  */
  assign n1145_o = x == 9'b000000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:43:13  */
  assign n1148_o = x == 9'b000000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:44:13  */
  assign n1151_o = x == 9'b000001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:45:13  */
  assign n1154_o = x == 9'b000001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:46:13  */
  assign n1157_o = x == 9'b000001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:47:13  */
  assign n1160_o = x == 9'b000001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:48:13  */
  assign n1163_o = x == 9'b000001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:49:13  */
  assign n1166_o = x == 9'b000001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:50:13  */
  assign n1169_o = x == 9'b000001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:51:13  */
  assign n1172_o = x == 9'b000001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:52:13  */
  assign n1175_o = x == 9'b000010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:53:13  */
  assign n1178_o = x == 9'b000010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:54:13  */
  assign n1181_o = x == 9'b000010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:55:13  */
  assign n1184_o = x == 9'b000010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:56:13  */
  assign n1187_o = x == 9'b000010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:57:13  */
  assign n1190_o = x == 9'b000010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:58:13  */
  assign n1193_o = x == 9'b000010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:59:13  */
  assign n1196_o = x == 9'b000010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:60:13  */
  assign n1199_o = x == 9'b000011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:61:13  */
  assign n1202_o = x == 9'b000011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:62:13  */
  assign n1205_o = x == 9'b000011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:63:13  */
  assign n1208_o = x == 9'b000011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:64:13  */
  assign n1211_o = x == 9'b000011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:65:13  */
  assign n1214_o = x == 9'b000011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:66:13  */
  assign n1217_o = x == 9'b000011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:67:13  */
  assign n1220_o = x == 9'b000011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:68:13  */
  assign n1223_o = x == 9'b000100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:69:13  */
  assign n1226_o = x == 9'b000100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:70:13  */
  assign n1229_o = x == 9'b000100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:71:13  */
  assign n1232_o = x == 9'b000100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:72:13  */
  assign n1235_o = x == 9'b000100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:73:13  */
  assign n1238_o = x == 9'b000100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:74:13  */
  assign n1241_o = x == 9'b000100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:75:13  */
  assign n1244_o = x == 9'b000100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:76:13  */
  assign n1247_o = x == 9'b000101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:77:13  */
  assign n1250_o = x == 9'b000101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:78:13  */
  assign n1253_o = x == 9'b000101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:79:13  */
  assign n1256_o = x == 9'b000101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:80:13  */
  assign n1259_o = x == 9'b000101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:81:13  */
  assign n1262_o = x == 9'b000101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:82:13  */
  assign n1265_o = x == 9'b000101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:83:13  */
  assign n1268_o = x == 9'b000101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:84:13  */
  assign n1271_o = x == 9'b000110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:85:13  */
  assign n1274_o = x == 9'b000110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:86:13  */
  assign n1277_o = x == 9'b000110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:87:13  */
  assign n1280_o = x == 9'b000110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:88:13  */
  assign n1283_o = x == 9'b000110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:89:13  */
  assign n1286_o = x == 9'b000110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:90:13  */
  assign n1289_o = x == 9'b000110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:91:13  */
  assign n1292_o = x == 9'b000110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:92:13  */
  assign n1295_o = x == 9'b000111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:93:13  */
  assign n1298_o = x == 9'b000111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:94:13  */
  assign n1301_o = x == 9'b000111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:95:13  */
  assign n1304_o = x == 9'b000111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:96:13  */
  assign n1307_o = x == 9'b000111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:97:13  */
  assign n1310_o = x == 9'b000111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:98:13  */
  assign n1313_o = x == 9'b000111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:99:13  */
  assign n1316_o = x == 9'b000111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:100:13  */
  assign n1319_o = x == 9'b001000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:101:13  */
  assign n1322_o = x == 9'b001000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:102:13  */
  assign n1325_o = x == 9'b001000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:103:13  */
  assign n1328_o = x == 9'b001000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:104:13  */
  assign n1331_o = x == 9'b001000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:105:13  */
  assign n1334_o = x == 9'b001000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:106:13  */
  assign n1337_o = x == 9'b001000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:107:13  */
  assign n1340_o = x == 9'b001000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:108:13  */
  assign n1343_o = x == 9'b001001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:109:13  */
  assign n1346_o = x == 9'b001001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:110:13  */
  assign n1349_o = x == 9'b001001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:111:13  */
  assign n1352_o = x == 9'b001001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:112:13  */
  assign n1355_o = x == 9'b001001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:113:13  */
  assign n1358_o = x == 9'b001001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:114:13  */
  assign n1361_o = x == 9'b001001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:115:13  */
  assign n1364_o = x == 9'b001001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:116:13  */
  assign n1367_o = x == 9'b001010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:117:13  */
  assign n1370_o = x == 9'b001010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:118:13  */
  assign n1373_o = x == 9'b001010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:119:13  */
  assign n1376_o = x == 9'b001010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:120:13  */
  assign n1379_o = x == 9'b001010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:121:13  */
  assign n1382_o = x == 9'b001010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:122:13  */
  assign n1385_o = x == 9'b001010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:123:13  */
  assign n1388_o = x == 9'b001010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:124:13  */
  assign n1391_o = x == 9'b001011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:125:13  */
  assign n1394_o = x == 9'b001011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:126:13  */
  assign n1397_o = x == 9'b001011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:127:13  */
  assign n1400_o = x == 9'b001011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:128:13  */
  assign n1403_o = x == 9'b001011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:129:13  */
  assign n1406_o = x == 9'b001011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:130:13  */
  assign n1409_o = x == 9'b001011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:131:13  */
  assign n1412_o = x == 9'b001011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:132:13  */
  assign n1415_o = x == 9'b001100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:133:13  */
  assign n1418_o = x == 9'b001100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:134:13  */
  assign n1421_o = x == 9'b001100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:135:13  */
  assign n1424_o = x == 9'b001100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:136:13  */
  assign n1427_o = x == 9'b001100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:137:13  */
  assign n1430_o = x == 9'b001100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:138:13  */
  assign n1433_o = x == 9'b001100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:139:13  */
  assign n1436_o = x == 9'b001100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:140:13  */
  assign n1439_o = x == 9'b001101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:141:13  */
  assign n1442_o = x == 9'b001101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:142:13  */
  assign n1445_o = x == 9'b001101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:143:13  */
  assign n1448_o = x == 9'b001101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:144:13  */
  assign n1451_o = x == 9'b001101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:145:13  */
  assign n1454_o = x == 9'b001101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:146:13  */
  assign n1457_o = x == 9'b001101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:147:13  */
  assign n1460_o = x == 9'b001101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:148:13  */
  assign n1463_o = x == 9'b001110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:149:13  */
  assign n1466_o = x == 9'b001110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:150:13  */
  assign n1469_o = x == 9'b001110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:151:13  */
  assign n1472_o = x == 9'b001110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:152:13  */
  assign n1475_o = x == 9'b001110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:153:13  */
  assign n1478_o = x == 9'b001110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:154:13  */
  assign n1481_o = x == 9'b001110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:155:13  */
  assign n1484_o = x == 9'b001110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:156:13  */
  assign n1487_o = x == 9'b001111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:157:13  */
  assign n1490_o = x == 9'b001111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:158:13  */
  assign n1493_o = x == 9'b001111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:159:13  */
  assign n1496_o = x == 9'b001111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:160:13  */
  assign n1499_o = x == 9'b001111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:161:13  */
  assign n1502_o = x == 9'b001111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:162:13  */
  assign n1505_o = x == 9'b001111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:163:13  */
  assign n1508_o = x == 9'b001111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:164:13  */
  assign n1511_o = x == 9'b010000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:165:13  */
  assign n1514_o = x == 9'b010000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:166:13  */
  assign n1517_o = x == 9'b010000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:167:13  */
  assign n1520_o = x == 9'b010000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:168:13  */
  assign n1523_o = x == 9'b010000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:169:13  */
  assign n1526_o = x == 9'b010000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:170:13  */
  assign n1529_o = x == 9'b010000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:171:13  */
  assign n1532_o = x == 9'b010000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:172:13  */
  assign n1535_o = x == 9'b010001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:173:13  */
  assign n1538_o = x == 9'b010001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:174:13  */
  assign n1541_o = x == 9'b010001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:175:13  */
  assign n1544_o = x == 9'b010001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:176:13  */
  assign n1547_o = x == 9'b010001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:177:13  */
  assign n1550_o = x == 9'b010001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:178:13  */
  assign n1553_o = x == 9'b010001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:179:13  */
  assign n1556_o = x == 9'b010001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:180:13  */
  assign n1559_o = x == 9'b010010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:181:13  */
  assign n1562_o = x == 9'b010010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:182:13  */
  assign n1565_o = x == 9'b010010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:183:13  */
  assign n1568_o = x == 9'b010010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:184:13  */
  assign n1571_o = x == 9'b010010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:185:13  */
  assign n1574_o = x == 9'b010010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:186:13  */
  assign n1577_o = x == 9'b010010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:187:13  */
  assign n1580_o = x == 9'b010010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:188:13  */
  assign n1583_o = x == 9'b010011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:189:13  */
  assign n1586_o = x == 9'b010011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:190:13  */
  assign n1589_o = x == 9'b010011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:191:13  */
  assign n1592_o = x == 9'b010011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:192:13  */
  assign n1595_o = x == 9'b010011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:193:13  */
  assign n1598_o = x == 9'b010011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:194:13  */
  assign n1601_o = x == 9'b010011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:195:13  */
  assign n1604_o = x == 9'b010011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:196:13  */
  assign n1607_o = x == 9'b010100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:197:13  */
  assign n1610_o = x == 9'b010100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:198:13  */
  assign n1613_o = x == 9'b010100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:199:13  */
  assign n1616_o = x == 9'b010100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:200:13  */
  assign n1619_o = x == 9'b010100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:201:13  */
  assign n1622_o = x == 9'b010100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:202:13  */
  assign n1625_o = x == 9'b010100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:203:13  */
  assign n1628_o = x == 9'b010100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:204:13  */
  assign n1631_o = x == 9'b010101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:205:13  */
  assign n1634_o = x == 9'b010101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:206:13  */
  assign n1637_o = x == 9'b010101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:207:13  */
  assign n1640_o = x == 9'b010101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:208:13  */
  assign n1643_o = x == 9'b010101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:209:13  */
  assign n1646_o = x == 9'b010101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:210:13  */
  assign n1649_o = x == 9'b010101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:211:13  */
  assign n1652_o = x == 9'b010101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:212:13  */
  assign n1655_o = x == 9'b010110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:213:13  */
  assign n1658_o = x == 9'b010110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:214:13  */
  assign n1661_o = x == 9'b010110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:215:13  */
  assign n1664_o = x == 9'b010110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:216:13  */
  assign n1667_o = x == 9'b010110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:217:13  */
  assign n1670_o = x == 9'b010110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:218:13  */
  assign n1673_o = x == 9'b010110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:219:13  */
  assign n1676_o = x == 9'b010110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:220:13  */
  assign n1679_o = x == 9'b010111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:221:13  */
  assign n1682_o = x == 9'b010111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:222:13  */
  assign n1685_o = x == 9'b010111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:223:13  */
  assign n1688_o = x == 9'b010111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:224:13  */
  assign n1691_o = x == 9'b010111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:225:13  */
  assign n1694_o = x == 9'b010111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:226:13  */
  assign n1697_o = x == 9'b010111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:227:13  */
  assign n1700_o = x == 9'b010111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:228:13  */
  assign n1703_o = x == 9'b011000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:229:13  */
  assign n1706_o = x == 9'b011000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:230:13  */
  assign n1709_o = x == 9'b011000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:231:13  */
  assign n1712_o = x == 9'b011000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:232:13  */
  assign n1715_o = x == 9'b011000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:233:13  */
  assign n1718_o = x == 9'b011000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:234:13  */
  assign n1721_o = x == 9'b011000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:235:13  */
  assign n1724_o = x == 9'b011000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:236:13  */
  assign n1727_o = x == 9'b011001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:237:13  */
  assign n1730_o = x == 9'b011001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:238:13  */
  assign n1733_o = x == 9'b011001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:239:13  */
  assign n1736_o = x == 9'b011001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:240:13  */
  assign n1739_o = x == 9'b011001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:241:13  */
  assign n1742_o = x == 9'b011001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:242:13  */
  assign n1745_o = x == 9'b011001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:243:13  */
  assign n1748_o = x == 9'b011001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:244:13  */
  assign n1751_o = x == 9'b011010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:245:13  */
  assign n1754_o = x == 9'b011010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:246:13  */
  assign n1757_o = x == 9'b011010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:247:13  */
  assign n1760_o = x == 9'b011010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:248:13  */
  assign n1763_o = x == 9'b011010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:249:13  */
  assign n1766_o = x == 9'b011010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:250:13  */
  assign n1769_o = x == 9'b011010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:251:13  */
  assign n1772_o = x == 9'b011010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:252:13  */
  assign n1775_o = x == 9'b011011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:253:13  */
  assign n1778_o = x == 9'b011011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:254:13  */
  assign n1781_o = x == 9'b011011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:255:13  */
  assign n1784_o = x == 9'b011011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:256:13  */
  assign n1787_o = x == 9'b011011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:257:13  */
  assign n1790_o = x == 9'b011011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:258:13  */
  assign n1793_o = x == 9'b011011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:259:13  */
  assign n1796_o = x == 9'b011011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:260:13  */
  assign n1799_o = x == 9'b011100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:261:13  */
  assign n1802_o = x == 9'b011100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:262:13  */
  assign n1805_o = x == 9'b011100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:263:13  */
  assign n1808_o = x == 9'b011100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:264:13  */
  assign n1811_o = x == 9'b011100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:265:13  */
  assign n1814_o = x == 9'b011100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:266:13  */
  assign n1817_o = x == 9'b011100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:267:13  */
  assign n1820_o = x == 9'b011100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:268:13  */
  assign n1823_o = x == 9'b011101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:269:13  */
  assign n1826_o = x == 9'b011101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:270:13  */
  assign n1829_o = x == 9'b011101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:271:13  */
  assign n1832_o = x == 9'b011101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:272:13  */
  assign n1835_o = x == 9'b011101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:273:13  */
  assign n1838_o = x == 9'b011101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:274:13  */
  assign n1841_o = x == 9'b011101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:275:13  */
  assign n1844_o = x == 9'b011101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:276:13  */
  assign n1847_o = x == 9'b011110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:277:13  */
  assign n1850_o = x == 9'b011110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:278:13  */
  assign n1853_o = x == 9'b011110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:279:13  */
  assign n1856_o = x == 9'b011110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:280:13  */
  assign n1859_o = x == 9'b011110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:281:13  */
  assign n1862_o = x == 9'b011110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:282:13  */
  assign n1865_o = x == 9'b011110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:283:13  */
  assign n1868_o = x == 9'b011110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:284:13  */
  assign n1871_o = x == 9'b011111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:285:13  */
  assign n1874_o = x == 9'b011111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:286:13  */
  assign n1877_o = x == 9'b011111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:287:13  */
  assign n1880_o = x == 9'b011111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:288:13  */
  assign n1883_o = x == 9'b011111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:289:13  */
  assign n1886_o = x == 9'b011111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:290:13  */
  assign n1889_o = x == 9'b011111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:291:13  */
  assign n1892_o = x == 9'b011111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:292:13  */
  assign n1895_o = x == 9'b100000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:293:13  */
  assign n1898_o = x == 9'b100000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:294:13  */
  assign n1901_o = x == 9'b100000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:295:13  */
  assign n1904_o = x == 9'b100000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:296:13  */
  assign n1907_o = x == 9'b100000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:297:13  */
  assign n1910_o = x == 9'b100000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:298:13  */
  assign n1913_o = x == 9'b100000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:299:13  */
  assign n1916_o = x == 9'b100000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:300:13  */
  assign n1919_o = x == 9'b100001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:301:13  */
  assign n1922_o = x == 9'b100001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:302:13  */
  assign n1925_o = x == 9'b100001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:303:13  */
  assign n1928_o = x == 9'b100001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:304:13  */
  assign n1931_o = x == 9'b100001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:305:13  */
  assign n1934_o = x == 9'b100001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:306:13  */
  assign n1937_o = x == 9'b100001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:307:13  */
  assign n1940_o = x == 9'b100001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:308:13  */
  assign n1943_o = x == 9'b100010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:309:13  */
  assign n1946_o = x == 9'b100010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:310:13  */
  assign n1949_o = x == 9'b100010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:311:13  */
  assign n1952_o = x == 9'b100010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:312:13  */
  assign n1955_o = x == 9'b100010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:313:13  */
  assign n1958_o = x == 9'b100010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:314:13  */
  assign n1961_o = x == 9'b100010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:315:13  */
  assign n1964_o = x == 9'b100010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:316:13  */
  assign n1967_o = x == 9'b100011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:317:13  */
  assign n1970_o = x == 9'b100011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:318:13  */
  assign n1973_o = x == 9'b100011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:319:13  */
  assign n1976_o = x == 9'b100011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:320:13  */
  assign n1979_o = x == 9'b100011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:321:13  */
  assign n1982_o = x == 9'b100011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:322:13  */
  assign n1985_o = x == 9'b100011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:323:13  */
  assign n1988_o = x == 9'b100011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:324:13  */
  assign n1991_o = x == 9'b100100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:325:13  */
  assign n1994_o = x == 9'b100100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:326:13  */
  assign n1997_o = x == 9'b100100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:327:13  */
  assign n2000_o = x == 9'b100100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:328:13  */
  assign n2003_o = x == 9'b100100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:329:13  */
  assign n2006_o = x == 9'b100100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:330:13  */
  assign n2009_o = x == 9'b100100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:331:13  */
  assign n2012_o = x == 9'b100100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:332:13  */
  assign n2015_o = x == 9'b100101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:333:13  */
  assign n2018_o = x == 9'b100101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:334:13  */
  assign n2021_o = x == 9'b100101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:335:13  */
  assign n2024_o = x == 9'b100101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:336:13  */
  assign n2027_o = x == 9'b100101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:337:13  */
  assign n2030_o = x == 9'b100101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:338:13  */
  assign n2033_o = x == 9'b100101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:339:13  */
  assign n2036_o = x == 9'b100101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:340:13  */
  assign n2039_o = x == 9'b100110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:341:13  */
  assign n2042_o = x == 9'b100110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:342:13  */
  assign n2045_o = x == 9'b100110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:343:13  */
  assign n2048_o = x == 9'b100110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:344:13  */
  assign n2051_o = x == 9'b100110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:345:13  */
  assign n2054_o = x == 9'b100110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:346:13  */
  assign n2057_o = x == 9'b100110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:347:13  */
  assign n2060_o = x == 9'b100110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:348:13  */
  assign n2063_o = x == 9'b100111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:349:13  */
  assign n2066_o = x == 9'b100111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:350:13  */
  assign n2069_o = x == 9'b100111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:351:13  */
  assign n2072_o = x == 9'b100111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:352:13  */
  assign n2075_o = x == 9'b100111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:353:13  */
  assign n2078_o = x == 9'b100111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:354:13  */
  assign n2081_o = x == 9'b100111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:355:13  */
  assign n2084_o = x == 9'b100111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:356:13  */
  assign n2087_o = x == 9'b101000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:357:13  */
  assign n2090_o = x == 9'b101000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:358:13  */
  assign n2093_o = x == 9'b101000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:359:13  */
  assign n2096_o = x == 9'b101000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:360:13  */
  assign n2099_o = x == 9'b101000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:361:13  */
  assign n2102_o = x == 9'b101000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:362:13  */
  assign n2105_o = x == 9'b101000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:363:13  */
  assign n2108_o = x == 9'b101000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:364:13  */
  assign n2111_o = x == 9'b101001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:365:13  */
  assign n2114_o = x == 9'b101001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:366:13  */
  assign n2117_o = x == 9'b101001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:367:13  */
  assign n2120_o = x == 9'b101001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:368:13  */
  assign n2123_o = x == 9'b101001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:369:13  */
  assign n2126_o = x == 9'b101001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:370:13  */
  assign n2129_o = x == 9'b101001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:371:13  */
  assign n2132_o = x == 9'b101001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:372:13  */
  assign n2135_o = x == 9'b101010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:373:13  */
  assign n2138_o = x == 9'b101010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:374:13  */
  assign n2141_o = x == 9'b101010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:375:13  */
  assign n2144_o = x == 9'b101010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:376:13  */
  assign n2147_o = x == 9'b101010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:377:13  */
  assign n2150_o = x == 9'b101010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:378:13  */
  assign n2153_o = x == 9'b101010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:379:13  */
  assign n2156_o = x == 9'b101010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:380:13  */
  assign n2159_o = x == 9'b101011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:381:13  */
  assign n2162_o = x == 9'b101011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:382:13  */
  assign n2165_o = x == 9'b101011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:383:13  */
  assign n2168_o = x == 9'b101011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:384:13  */
  assign n2171_o = x == 9'b101011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:385:13  */
  assign n2174_o = x == 9'b101011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:386:13  */
  assign n2177_o = x == 9'b101011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:387:13  */
  assign n2180_o = x == 9'b101011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:388:13  */
  assign n2183_o = x == 9'b101100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:389:13  */
  assign n2186_o = x == 9'b101100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:390:13  */
  assign n2189_o = x == 9'b101100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:391:13  */
  assign n2192_o = x == 9'b101100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:392:13  */
  assign n2195_o = x == 9'b101100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:393:13  */
  assign n2198_o = x == 9'b101100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:394:13  */
  assign n2201_o = x == 9'b101100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:395:13  */
  assign n2204_o = x == 9'b101100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:396:13  */
  assign n2207_o = x == 9'b101101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:397:13  */
  assign n2210_o = x == 9'b101101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:398:13  */
  assign n2213_o = x == 9'b101101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:399:13  */
  assign n2216_o = x == 9'b101101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:400:13  */
  assign n2219_o = x == 9'b101101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:401:13  */
  assign n2222_o = x == 9'b101101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:402:13  */
  assign n2225_o = x == 9'b101101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:403:13  */
  assign n2228_o = x == 9'b101101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:404:13  */
  assign n2231_o = x == 9'b101110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:405:13  */
  assign n2234_o = x == 9'b101110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:406:13  */
  assign n2237_o = x == 9'b101110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:407:13  */
  assign n2240_o = x == 9'b101110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:408:13  */
  assign n2243_o = x == 9'b101110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:409:13  */
  assign n2246_o = x == 9'b101110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:410:13  */
  assign n2249_o = x == 9'b101110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:411:13  */
  assign n2252_o = x == 9'b101110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:412:13  */
  assign n2255_o = x == 9'b101111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:413:13  */
  assign n2258_o = x == 9'b101111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:414:13  */
  assign n2261_o = x == 9'b101111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:415:13  */
  assign n2264_o = x == 9'b101111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:416:13  */
  assign n2267_o = x == 9'b101111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:417:13  */
  assign n2270_o = x == 9'b101111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:418:13  */
  assign n2273_o = x == 9'b101111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:419:13  */
  assign n2276_o = x == 9'b101111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:420:13  */
  assign n2279_o = x == 9'b110000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:421:13  */
  assign n2282_o = x == 9'b110000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:422:13  */
  assign n2285_o = x == 9'b110000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:423:13  */
  assign n2288_o = x == 9'b110000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:424:13  */
  assign n2291_o = x == 9'b110000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:425:13  */
  assign n2294_o = x == 9'b110000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:426:13  */
  assign n2297_o = x == 9'b110000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:427:13  */
  assign n2300_o = x == 9'b110000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:428:13  */
  assign n2303_o = x == 9'b110001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:429:13  */
  assign n2306_o = x == 9'b110001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:430:13  */
  assign n2309_o = x == 9'b110001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:431:13  */
  assign n2312_o = x == 9'b110001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:432:13  */
  assign n2315_o = x == 9'b110001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:433:13  */
  assign n2318_o = x == 9'b110001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:434:13  */
  assign n2321_o = x == 9'b110001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:435:13  */
  assign n2324_o = x == 9'b110001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:436:13  */
  assign n2327_o = x == 9'b110010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:437:13  */
  assign n2330_o = x == 9'b110010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:438:13  */
  assign n2333_o = x == 9'b110010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:439:13  */
  assign n2336_o = x == 9'b110010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:440:13  */
  assign n2339_o = x == 9'b110010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:441:13  */
  assign n2342_o = x == 9'b110010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:442:13  */
  assign n2345_o = x == 9'b110010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:443:13  */
  assign n2348_o = x == 9'b110010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:444:13  */
  assign n2351_o = x == 9'b110011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:445:13  */
  assign n2354_o = x == 9'b110011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:446:13  */
  assign n2357_o = x == 9'b110011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:447:13  */
  assign n2360_o = x == 9'b110011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:448:13  */
  assign n2363_o = x == 9'b110011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:449:13  */
  assign n2366_o = x == 9'b110011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:450:13  */
  assign n2369_o = x == 9'b110011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:451:13  */
  assign n2372_o = x == 9'b110011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:452:13  */
  assign n2375_o = x == 9'b110100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:453:13  */
  assign n2378_o = x == 9'b110100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:454:13  */
  assign n2381_o = x == 9'b110100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:455:13  */
  assign n2384_o = x == 9'b110100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:456:13  */
  assign n2387_o = x == 9'b110100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:457:13  */
  assign n2390_o = x == 9'b110100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:458:13  */
  assign n2393_o = x == 9'b110100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:459:13  */
  assign n2396_o = x == 9'b110100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:460:13  */
  assign n2399_o = x == 9'b110101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:461:13  */
  assign n2402_o = x == 9'b110101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:462:13  */
  assign n2405_o = x == 9'b110101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:463:13  */
  assign n2408_o = x == 9'b110101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:464:13  */
  assign n2411_o = x == 9'b110101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:465:13  */
  assign n2414_o = x == 9'b110101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:466:13  */
  assign n2417_o = x == 9'b110101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:467:13  */
  assign n2420_o = x == 9'b110101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:468:13  */
  assign n2423_o = x == 9'b110110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:469:13  */
  assign n2426_o = x == 9'b110110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:470:13  */
  assign n2429_o = x == 9'b110110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:471:13  */
  assign n2432_o = x == 9'b110110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:472:13  */
  assign n2435_o = x == 9'b110110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:473:13  */
  assign n2438_o = x == 9'b110110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:474:13  */
  assign n2441_o = x == 9'b110110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:475:13  */
  assign n2444_o = x == 9'b110110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:476:13  */
  assign n2447_o = x == 9'b110111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:477:13  */
  assign n2450_o = x == 9'b110111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:478:13  */
  assign n2453_o = x == 9'b110111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:479:13  */
  assign n2456_o = x == 9'b110111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:480:13  */
  assign n2459_o = x == 9'b110111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:481:13  */
  assign n2462_o = x == 9'b110111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:482:13  */
  assign n2465_o = x == 9'b110111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:483:13  */
  assign n2468_o = x == 9'b110111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:484:13  */
  assign n2471_o = x == 9'b111000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:485:13  */
  assign n2474_o = x == 9'b111000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:486:13  */
  assign n2477_o = x == 9'b111000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:487:13  */
  assign n2480_o = x == 9'b111000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:488:13  */
  assign n2483_o = x == 9'b111000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:489:13  */
  assign n2486_o = x == 9'b111000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:490:13  */
  assign n2489_o = x == 9'b111000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:491:13  */
  assign n2492_o = x == 9'b111000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:492:13  */
  assign n2495_o = x == 9'b111001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:493:13  */
  assign n2498_o = x == 9'b111001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:494:13  */
  assign n2501_o = x == 9'b111001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:495:13  */
  assign n2504_o = x == 9'b111001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:496:13  */
  assign n2507_o = x == 9'b111001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:497:13  */
  assign n2510_o = x == 9'b111001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:498:13  */
  assign n2513_o = x == 9'b111001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:499:13  */
  assign n2516_o = x == 9'b111001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:500:13  */
  assign n2519_o = x == 9'b111010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:501:13  */
  assign n2522_o = x == 9'b111010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:502:13  */
  assign n2525_o = x == 9'b111010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:503:13  */
  assign n2528_o = x == 9'b111010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:504:13  */
  assign n2531_o = x == 9'b111010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:505:13  */
  assign n2534_o = x == 9'b111010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:506:13  */
  assign n2537_o = x == 9'b111010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:507:13  */
  assign n2540_o = x == 9'b111010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:508:13  */
  assign n2543_o = x == 9'b111011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:509:13  */
  assign n2546_o = x == 9'b111011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:510:13  */
  assign n2549_o = x == 9'b111011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:511:13  */
  assign n2552_o = x == 9'b111011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:512:13  */
  assign n2555_o = x == 9'b111011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:513:13  */
  assign n2558_o = x == 9'b111011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:514:13  */
  assign n2561_o = x == 9'b111011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:515:13  */
  assign n2564_o = x == 9'b111011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:516:13  */
  assign n2567_o = x == 9'b111100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:517:13  */
  assign n2570_o = x == 9'b111100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:518:13  */
  assign n2573_o = x == 9'b111100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:519:13  */
  assign n2576_o = x == 9'b111100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:520:13  */
  assign n2579_o = x == 9'b111100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:521:13  */
  assign n2582_o = x == 9'b111100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:522:13  */
  assign n2585_o = x == 9'b111100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:523:13  */
  assign n2588_o = x == 9'b111100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:524:13  */
  assign n2591_o = x == 9'b111101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:525:13  */
  assign n2594_o = x == 9'b111101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:526:13  */
  assign n2597_o = x == 9'b111101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:527:13  */
  assign n2600_o = x == 9'b111101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:528:13  */
  assign n2603_o = x == 9'b111101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:529:13  */
  assign n2606_o = x == 9'b111101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:530:13  */
  assign n2609_o = x == 9'b111101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:531:13  */
  assign n2612_o = x == 9'b111101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:532:13  */
  assign n2615_o = x == 9'b111110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:533:13  */
  assign n2618_o = x == 9'b111110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:534:13  */
  assign n2621_o = x == 9'b111110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:535:13  */
  assign n2624_o = x == 9'b111110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:536:13  */
  assign n2627_o = x == 9'b111110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:537:13  */
  assign n2630_o = x == 9'b111110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:538:13  */
  assign n2633_o = x == 9'b111110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:539:13  */
  assign n2636_o = x == 9'b111110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:540:13  */
  assign n2639_o = x == 9'b111111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:541:13  */
  assign n2642_o = x == 9'b111111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:542:13  */
  assign n2645_o = x == 9'b111111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:543:13  */
  assign n2648_o = x == 9'b111111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:544:13  */
  assign n2651_o = x == 9'b111111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:545:13  */
  assign n2654_o = x == 9'b111111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:546:13  */
  assign n2657_o = x == 9'b111111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:547:13  */
  assign n2660_o = x == 9'b111111111;
  assign n2662_o = {n2660_o, n2657_o, n2654_o, n2651_o, n2648_o, n2645_o, n2642_o, n2639_o, n2636_o, n2633_o, n2630_o, n2627_o, n2624_o, n2621_o, n2618_o, n2615_o, n2612_o, n2609_o, n2606_o, n2603_o, n2600_o, n2597_o, n2594_o, n2591_o, n2588_o, n2585_o, n2582_o, n2579_o, n2576_o, n2573_o, n2570_o, n2567_o, n2564_o, n2561_o, n2558_o, n2555_o, n2552_o, n2549_o, n2546_o, n2543_o, n2540_o, n2537_o, n2534_o, n2531_o, n2528_o, n2525_o, n2522_o, n2519_o, n2516_o, n2513_o, n2510_o, n2507_o, n2504_o, n2501_o, n2498_o, n2495_o, n2492_o, n2489_o, n2486_o, n2483_o, n2480_o, n2477_o, n2474_o, n2471_o, n2468_o, n2465_o, n2462_o, n2459_o, n2456_o, n2453_o, n2450_o, n2447_o, n2444_o, n2441_o, n2438_o, n2435_o, n2432_o, n2429_o, n2426_o, n2423_o, n2420_o, n2417_o, n2414_o, n2411_o, n2408_o, n2405_o, n2402_o, n2399_o, n2396_o, n2393_o, n2390_o, n2387_o, n2384_o, n2381_o, n2378_o, n2375_o, n2372_o, n2369_o, n2366_o, n2363_o, n2360_o, n2357_o, n2354_o, n2351_o, n2348_o, n2345_o, n2342_o, n2339_o, n2336_o, n2333_o, n2330_o, n2327_o, n2324_o, n2321_o, n2318_o, n2315_o, n2312_o, n2309_o, n2306_o, n2303_o, n2300_o, n2297_o, n2294_o, n2291_o, n2288_o, n2285_o, n2282_o, n2279_o, n2276_o, n2273_o, n2270_o, n2267_o, n2264_o, n2261_o, n2258_o, n2255_o, n2252_o, n2249_o, n2246_o, n2243_o, n2240_o, n2237_o, n2234_o, n2231_o, n2228_o, n2225_o, n2222_o, n2219_o, n2216_o, n2213_o, n2210_o, n2207_o, n2204_o, n2201_o, n2198_o, n2195_o, n2192_o, n2189_o, n2186_o, n2183_o, n2180_o, n2177_o, n2174_o, n2171_o, n2168_o, n2165_o, n2162_o, n2159_o, n2156_o, n2153_o, n2150_o, n2147_o, n2144_o, n2141_o, n2138_o, n2135_o, n2132_o, n2129_o, n2126_o, n2123_o, n2120_o, n2117_o, n2114_o, n2111_o, n2108_o, n2105_o, n2102_o, n2099_o, n2096_o, n2093_o, n2090_o, n2087_o, n2084_o, n2081_o, n2078_o, n2075_o, n2072_o, n2069_o, n2066_o, n2063_o, n2060_o, n2057_o, n2054_o, n2051_o, n2048_o, n2045_o, n2042_o, n2039_o, n2036_o, n2033_o, n2030_o, n2027_o, n2024_o, n2021_o, n2018_o, n2015_o, n2012_o, n2009_o, n2006_o, n2003_o, n2000_o, n1997_o, n1994_o, n1991_o, n1988_o, n1985_o, n1982_o, n1979_o, n1976_o, n1973_o, n1970_o, n1967_o, n1964_o, n1961_o, n1958_o, n1955_o, n1952_o, n1949_o, n1946_o, n1943_o, n1940_o, n1937_o, n1934_o, n1931_o, n1928_o, n1925_o, n1922_o, n1919_o, n1916_o, n1913_o, n1910_o, n1907_o, n1904_o, n1901_o, n1898_o, n1895_o, n1892_o, n1889_o, n1886_o, n1883_o, n1880_o, n1877_o, n1874_o, n1871_o, n1868_o, n1865_o, n1862_o, n1859_o, n1856_o, n1853_o, n1850_o, n1847_o, n1844_o, n1841_o, n1838_o, n1835_o, n1832_o, n1829_o, n1826_o, n1823_o, n1820_o, n1817_o, n1814_o, n1811_o, n1808_o, n1805_o, n1802_o, n1799_o, n1796_o, n1793_o, n1790_o, n1787_o, n1784_o, n1781_o, n1778_o, n1775_o, n1772_o, n1769_o, n1766_o, n1763_o, n1760_o, n1757_o, n1754_o, n1751_o, n1748_o, n1745_o, n1742_o, n1739_o, n1736_o, n1733_o, n1730_o, n1727_o, n1724_o, n1721_o, n1718_o, n1715_o, n1712_o, n1709_o, n1706_o, n1703_o, n1700_o, n1697_o, n1694_o, n1691_o, n1688_o, n1685_o, n1682_o, n1679_o, n1676_o, n1673_o, n1670_o, n1667_o, n1664_o, n1661_o, n1658_o, n1655_o, n1652_o, n1649_o, n1646_o, n1643_o, n1640_o, n1637_o, n1634_o, n1631_o, n1628_o, n1625_o, n1622_o, n1619_o, n1616_o, n1613_o, n1610_o, n1607_o, n1604_o, n1601_o, n1598_o, n1595_o, n1592_o, n1589_o, n1586_o, n1583_o, n1580_o, n1577_o, n1574_o, n1571_o, n1568_o, n1565_o, n1562_o, n1559_o, n1556_o, n1553_o, n1550_o, n1547_o, n1544_o, n1541_o, n1538_o, n1535_o, n1532_o, n1529_o, n1526_o, n1523_o, n1520_o, n1517_o, n1514_o, n1511_o, n1508_o, n1505_o, n1502_o, n1499_o, n1496_o, n1493_o, n1490_o, n1487_o, n1484_o, n1481_o, n1478_o, n1475_o, n1472_o, n1469_o, n1466_o, n1463_o, n1460_o, n1457_o, n1454_o, n1451_o, n1448_o, n1445_o, n1442_o, n1439_o, n1436_o, n1433_o, n1430_o, n1427_o, n1424_o, n1421_o, n1418_o, n1415_o, n1412_o, n1409_o, n1406_o, n1403_o, n1400_o, n1397_o, n1394_o, n1391_o, n1388_o, n1385_o, n1382_o, n1379_o, n1376_o, n1373_o, n1370_o, n1367_o, n1364_o, n1361_o, n1358_o, n1355_o, n1352_o, n1349_o, n1346_o, n1343_o, n1340_o, n1337_o, n1334_o, n1331_o, n1328_o, n1325_o, n1322_o, n1319_o, n1316_o, n1313_o, n1310_o, n1307_o, n1304_o, n1301_o, n1298_o, n1295_o, n1292_o, n1289_o, n1286_o, n1283_o, n1280_o, n1277_o, n1274_o, n1271_o, n1268_o, n1265_o, n1262_o, n1259_o, n1256_o, n1253_o, n1250_o, n1247_o, n1244_o, n1241_o, n1238_o, n1235_o, n1232_o, n1229_o, n1226_o, n1223_o, n1220_o, n1217_o, n1214_o, n1211_o, n1208_o, n1205_o, n1202_o, n1199_o, n1196_o, n1193_o, n1190_o, n1187_o, n1184_o, n1181_o, n1178_o, n1175_o, n1172_o, n1169_o, n1166_o, n1163_o, n1160_o, n1157_o, n1154_o, n1151_o, n1148_o, n1145_o, n1142_o, n1139_o, n1136_o, n1133_o, n1130_o, n1127_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:35:4  */
  always @*
    case (n2662_o)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2663_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2663_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2663_o = 3'b000;
      default: n2663_o = 3'bXXX;
    endcase
endmodule

module fdiv #(parameter ID = 1)
  (input  clk,
   input  [33:0] X,
   input  [33:0] Y,
   output [33:0] R);
  wire [23:0] fx;
  wire [23:0] fy;
  wire [9:0] expr0;
  wire [9:0] expr0_d1;
  wire [9:0] expr0_d2;
  wire [9:0] expr0_d3;
  wire [9:0] expr0_d4;
  wire [9:0] expr0_d5;
  wire [9:0] expr0_d6;
  wire [9:0] expr0_d7;
  wire [9:0] expr0_d8;
  wire [9:0] expr0_d9;
  wire [9:0] expr0_d10;
  wire [9:0] expr0_d11;
  wire [9:0] expr0_d12;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire sr_d7;
  wire sr_d8;
  wire sr_d9;
  wire sr_d10;
  wire sr_d11;
  wire sr_d12;
  wire [3:0] exnxy;
  wire [1:0] exnr0;
  wire [1:0] exnr0_d1;
  wire [1:0] exnr0_d2;
  wire [1:0] exnr0_d3;
  wire [1:0] exnr0_d4;
  wire [1:0] exnr0_d5;
  wire [1:0] exnr0_d6;
  wire [1:0] exnr0_d7;
  wire [1:0] exnr0_d8;
  wire [1:0] exnr0_d9;
  wire [1:0] exnr0_d10;
  wire [1:0] exnr0_d11;
  wire [1:0] exnr0_d12;
  wire [23:0] d;
  wire [23:0] d_d1;
  wire [23:0] d_d2;
  wire [23:0] d_d3;
  wire [23:0] d_d4;
  wire [23:0] d_d5;
  wire [23:0] d_d6;
  wire [23:0] d_d7;
  wire [23:0] d_d8;
  wire [23:0] d_d9;
  wire [23:0] d_d10;
  wire [23:0] d_d11;
  wire [24:0] psx;
  wire [26:0] betaw14;
  wire [8:0] sel14;
  wire [2:0] q14;
  wire [2:0] q14_copy5;
  wire [26:0] absq14d;
  wire [26:0] w13;
  wire [26:0] betaw13;
  wire [26:0] betaw13_d1;
  wire [8:0] sel13;
  wire [2:0] q13;
  wire [2:0] q13_copy6;
  wire [2:0] q13_copy6_d1;
  wire [26:0] absq13d;
  wire [26:0] w12;
  wire [26:0] betaw12;
  wire [26:0] betaw12_d1;
  wire [8:0] sel12;
  wire [2:0] q12;
  wire [2:0] q12_copy7;
  wire [2:0] q12_copy7_d1;
  wire [26:0] absq12d;
  wire [26:0] w11;
  wire [26:0] betaw11;
  wire [26:0] betaw11_d1;
  wire [8:0] sel11;
  wire [2:0] q11;
  wire [2:0] q11_copy8;
  wire [2:0] q11_copy8_d1;
  wire [26:0] absq11d;
  wire [26:0] w10;
  wire [26:0] betaw10;
  wire [26:0] betaw10_d1;
  wire [8:0] sel10;
  wire [2:0] q10;
  wire [2:0] q10_d1;
  wire [2:0] q10_copy9;
  wire [26:0] absq10d;
  wire [26:0] absq10d_d1;
  wire [26:0] w9;
  wire [26:0] betaw9;
  wire [26:0] betaw9_d1;
  wire [8:0] sel9;
  wire [2:0] q9;
  wire [2:0] q9_d1;
  wire [2:0] q9_copy10;
  wire [26:0] absq9d;
  wire [26:0] absq9d_d1;
  wire [26:0] w8;
  wire [26:0] betaw8;
  wire [26:0] betaw8_d1;
  wire [8:0] sel8;
  wire [2:0] q8;
  wire [2:0] q8_d1;
  wire [2:0] q8_copy11;
  wire [26:0] absq8d;
  wire [26:0] absq8d_d1;
  wire [26:0] w7;
  wire [26:0] betaw7;
  wire [8:0] sel7;
  wire [2:0] q7;
  wire [2:0] q7_copy12;
  wire [26:0] absq7d;
  wire [26:0] w6;
  wire [26:0] betaw6;
  wire [26:0] betaw6_d1;
  wire [8:0] sel6;
  wire [2:0] q6;
  wire [2:0] q6_copy13;
  wire [2:0] q6_copy13_d1;
  wire [26:0] absq6d;
  wire [26:0] w5;
  wire [26:0] betaw5;
  wire [26:0] betaw5_d1;
  wire [8:0] sel5;
  wire [2:0] q5;
  wire [2:0] q5_copy14;
  wire [2:0] q5_copy14_d1;
  wire [26:0] absq5d;
  wire [26:0] w4;
  wire [26:0] betaw4;
  wire [26:0] betaw4_d1;
  wire [8:0] sel4;
  wire [2:0] q4;
  wire [2:0] q4_copy15;
  wire [2:0] q4_copy15_d1;
  wire [26:0] absq4d;
  wire [26:0] w3;
  wire [26:0] betaw3;
  wire [26:0] betaw3_d1;
  wire [8:0] sel3;
  wire [2:0] q3;
  wire [2:0] q3_copy16;
  wire [2:0] q3_copy16_d1;
  wire [26:0] absq3d;
  wire [26:0] w2;
  wire [26:0] betaw2;
  wire [26:0] betaw2_d1;
  wire [8:0] sel2;
  wire [2:0] q2;
  wire [2:0] q2_d1;
  wire [2:0] q2_copy17;
  wire [26:0] absq2d;
  wire [26:0] absq2d_d1;
  wire [26:0] w1;
  wire [26:0] betaw1;
  wire [26:0] betaw1_d1;
  wire [8:0] sel1;
  wire [2:0] q1;
  wire [2:0] q1_d1;
  wire [2:0] q1_copy18;
  wire [26:0] absq1d;
  wire [26:0] absq1d_d1;
  wire [26:0] w0;
  wire [24:0] wfinal;
  wire qm0;
  wire [1:0] qp14;
  wire [1:0] qp14_d1;
  wire [1:0] qp14_d2;
  wire [1:0] qp14_d3;
  wire [1:0] qp14_d4;
  wire [1:0] qp14_d5;
  wire [1:0] qp14_d6;
  wire [1:0] qp14_d7;
  wire [1:0] qp14_d8;
  wire [1:0] qp14_d9;
  wire [1:0] qp14_d10;
  wire [1:0] qp14_d11;
  wire [1:0] qm14;
  wire [1:0] qm14_d1;
  wire [1:0] qm14_d2;
  wire [1:0] qm14_d3;
  wire [1:0] qm14_d4;
  wire [1:0] qm14_d5;
  wire [1:0] qm14_d6;
  wire [1:0] qm14_d7;
  wire [1:0] qm14_d8;
  wire [1:0] qm14_d9;
  wire [1:0] qm14_d10;
  wire [1:0] qm14_d11;
  wire [1:0] qm14_d12;
  wire [1:0] qp13;
  wire [1:0] qp13_d1;
  wire [1:0] qp13_d2;
  wire [1:0] qp13_d3;
  wire [1:0] qp13_d4;
  wire [1:0] qp13_d5;
  wire [1:0] qp13_d6;
  wire [1:0] qp13_d7;
  wire [1:0] qp13_d8;
  wire [1:0] qp13_d9;
  wire [1:0] qp13_d10;
  wire [1:0] qm13;
  wire [1:0] qm13_d1;
  wire [1:0] qm13_d2;
  wire [1:0] qm13_d3;
  wire [1:0] qm13_d4;
  wire [1:0] qm13_d5;
  wire [1:0] qm13_d6;
  wire [1:0] qm13_d7;
  wire [1:0] qm13_d8;
  wire [1:0] qm13_d9;
  wire [1:0] qm13_d10;
  wire [1:0] qm13_d11;
  wire [1:0] qp12;
  wire [1:0] qp12_d1;
  wire [1:0] qp12_d2;
  wire [1:0] qp12_d3;
  wire [1:0] qp12_d4;
  wire [1:0] qp12_d5;
  wire [1:0] qp12_d6;
  wire [1:0] qp12_d7;
  wire [1:0] qp12_d8;
  wire [1:0] qp12_d9;
  wire [1:0] qm12;
  wire [1:0] qm12_d1;
  wire [1:0] qm12_d2;
  wire [1:0] qm12_d3;
  wire [1:0] qm12_d4;
  wire [1:0] qm12_d5;
  wire [1:0] qm12_d6;
  wire [1:0] qm12_d7;
  wire [1:0] qm12_d8;
  wire [1:0] qm12_d9;
  wire [1:0] qm12_d10;
  wire [1:0] qp11;
  wire [1:0] qp11_d1;
  wire [1:0] qp11_d2;
  wire [1:0] qp11_d3;
  wire [1:0] qp11_d4;
  wire [1:0] qp11_d5;
  wire [1:0] qp11_d6;
  wire [1:0] qp11_d7;
  wire [1:0] qp11_d8;
  wire [1:0] qm11;
  wire [1:0] qm11_d1;
  wire [1:0] qm11_d2;
  wire [1:0] qm11_d3;
  wire [1:0] qm11_d4;
  wire [1:0] qm11_d5;
  wire [1:0] qm11_d6;
  wire [1:0] qm11_d7;
  wire [1:0] qm11_d8;
  wire [1:0] qm11_d9;
  wire [1:0] qp10;
  wire [1:0] qp10_d1;
  wire [1:0] qp10_d2;
  wire [1:0] qp10_d3;
  wire [1:0] qp10_d4;
  wire [1:0] qp10_d5;
  wire [1:0] qp10_d6;
  wire [1:0] qp10_d7;
  wire [1:0] qp10_d8;
  wire [1:0] qm10;
  wire [1:0] qm10_d1;
  wire [1:0] qm10_d2;
  wire [1:0] qm10_d3;
  wire [1:0] qm10_d4;
  wire [1:0] qm10_d5;
  wire [1:0] qm10_d6;
  wire [1:0] qm10_d7;
  wire [1:0] qm10_d8;
  wire [1:0] qm10_d9;
  wire [1:0] qp9;
  wire [1:0] qp9_d1;
  wire [1:0] qp9_d2;
  wire [1:0] qp9_d3;
  wire [1:0] qp9_d4;
  wire [1:0] qp9_d5;
  wire [1:0] qp9_d6;
  wire [1:0] qp9_d7;
  wire [1:0] qm9;
  wire [1:0] qm9_d1;
  wire [1:0] qm9_d2;
  wire [1:0] qm9_d3;
  wire [1:0] qm9_d4;
  wire [1:0] qm9_d5;
  wire [1:0] qm9_d6;
  wire [1:0] qm9_d7;
  wire [1:0] qm9_d8;
  wire [1:0] qp8;
  wire [1:0] qp8_d1;
  wire [1:0] qp8_d2;
  wire [1:0] qp8_d3;
  wire [1:0] qp8_d4;
  wire [1:0] qp8_d5;
  wire [1:0] qp8_d6;
  wire [1:0] qm8;
  wire [1:0] qm8_d1;
  wire [1:0] qm8_d2;
  wire [1:0] qm8_d3;
  wire [1:0] qm8_d4;
  wire [1:0] qm8_d5;
  wire [1:0] qm8_d6;
  wire [1:0] qm8_d7;
  wire [1:0] qp7;
  wire [1:0] qp7_d1;
  wire [1:0] qp7_d2;
  wire [1:0] qp7_d3;
  wire [1:0] qp7_d4;
  wire [1:0] qp7_d5;
  wire [1:0] qm7;
  wire [1:0] qm7_d1;
  wire [1:0] qm7_d2;
  wire [1:0] qm7_d3;
  wire [1:0] qm7_d4;
  wire [1:0] qm7_d5;
  wire [1:0] qm7_d6;
  wire [1:0] qp6;
  wire [1:0] qp6_d1;
  wire [1:0] qp6_d2;
  wire [1:0] qp6_d3;
  wire [1:0] qp6_d4;
  wire [1:0] qm6;
  wire [1:0] qm6_d1;
  wire [1:0] qm6_d2;
  wire [1:0] qm6_d3;
  wire [1:0] qm6_d4;
  wire [1:0] qm6_d5;
  wire [1:0] qp5;
  wire [1:0] qp5_d1;
  wire [1:0] qp5_d2;
  wire [1:0] qp5_d3;
  wire [1:0] qm5;
  wire [1:0] qm5_d1;
  wire [1:0] qm5_d2;
  wire [1:0] qm5_d3;
  wire [1:0] qm5_d4;
  wire [1:0] qp4;
  wire [1:0] qp4_d1;
  wire [1:0] qp4_d2;
  wire [1:0] qm4;
  wire [1:0] qm4_d1;
  wire [1:0] qm4_d2;
  wire [1:0] qm4_d3;
  wire [1:0] qp3;
  wire [1:0] qp3_d1;
  wire [1:0] qm3;
  wire [1:0] qm3_d1;
  wire [1:0] qm3_d2;
  wire [1:0] qp2;
  wire [1:0] qp2_d1;
  wire [1:0] qm2;
  wire [1:0] qm2_d1;
  wire [1:0] qm2_d2;
  wire [1:0] qp1;
  wire [1:0] qm1;
  wire [1:0] qm1_d1;
  wire [27:0] qp;
  wire [27:0] qp_d1;
  wire [27:0] qm;
  wire [27:0] quotient;
  wire [25:0] mr;
  wire [23:0] frnorm;
  wire round;
  wire [9:0] expr1;
  wire [32:0] expfrac;
  wire [32:0] expfracr;
  wire [1:0] exnr;
  wire [1:0] exnrfinal;
  wire [22:0] n246_o;
  wire [23:0] n248_o;
  wire [22:0] n249_o;
  wire [23:0] n251_o;
  wire [7:0] n252_o;
  wire [9:0] n254_o;
  wire [7:0] n255_o;
  wire [9:0] n257_o;
  wire [9:0] n258_o;
  wire n259_o;
  wire n260_o;
  wire n261_o;
  wire [1:0] n262_o;
  wire [1:0] n263_o;
  wire [3:0] n264_o;
  wire n267_o;
  wire n270_o;
  wire n272_o;
  wire n273_o;
  wire n275_o;
  wire n276_o;
  wire n279_o;
  wire n281_o;
  wire n282_o;
  wire n284_o;
  wire n285_o;
  wire [2:0] n287_o;
  reg [1:0] n288_o;
  wire [24:0] n290_o;
  wire [26:0] n292_o;
  wire [5:0] n293_o;
  wire [2:0] n294_o;
  wire [8:0] n295_o;
  wire [2:0] selfunctiontable14_n296;
  wire [2:0] selfunctiontable14_y;
  wire [26:0] n300_o;
  wire n302_o;
  wire n304_o;
  wire n305_o;
  wire [25:0] n307_o;
  wire [26:0] n309_o;
  wire n311_o;
  wire n313_o;
  wire n314_o;
  wire [1:0] n316_o;
  reg [26:0] n317_o;
  wire n318_o;
  wire [26:0] n319_o;
  wire n321_o;
  wire [26:0] n322_o;
  reg [26:0] n323_o;
  wire [24:0] n324_o;
  wire [26:0] n326_o;
  wire [5:0] n327_o;
  wire [2:0] n328_o;
  wire [8:0] n329_o;
  wire [2:0] selfunctiontable13_n330;
  wire [2:0] selfunctiontable13_y;
  wire [26:0] n334_o;
  wire n336_o;
  wire n338_o;
  wire n339_o;
  wire [25:0] n341_o;
  wire [26:0] n343_o;
  wire n345_o;
  wire n347_o;
  wire n348_o;
  wire [1:0] n350_o;
  reg [26:0] n351_o;
  wire n352_o;
  wire [26:0] n353_o;
  wire n355_o;
  wire [26:0] n356_o;
  reg [26:0] n357_o;
  wire [24:0] n358_o;
  wire [26:0] n360_o;
  wire [5:0] n361_o;
  wire [2:0] n362_o;
  wire [8:0] n363_o;
  wire [2:0] selfunctiontable12_n364;
  wire [2:0] selfunctiontable12_y;
  wire [26:0] n368_o;
  wire n370_o;
  wire n372_o;
  wire n373_o;
  wire [25:0] n375_o;
  wire [26:0] n377_o;
  wire n379_o;
  wire n381_o;
  wire n382_o;
  wire [1:0] n384_o;
  reg [26:0] n385_o;
  wire n386_o;
  wire [26:0] n387_o;
  wire n389_o;
  wire [26:0] n390_o;
  reg [26:0] n391_o;
  wire [24:0] n392_o;
  wire [26:0] n394_o;
  wire [5:0] n395_o;
  wire [2:0] n396_o;
  wire [8:0] n397_o;
  wire [2:0] selfunctiontable11_n398;
  wire [2:0] selfunctiontable11_y;
  wire [26:0] n402_o;
  wire n404_o;
  wire n406_o;
  wire n407_o;
  wire [25:0] n409_o;
  wire [26:0] n411_o;
  wire n413_o;
  wire n415_o;
  wire n416_o;
  wire [1:0] n418_o;
  reg [26:0] n419_o;
  wire n420_o;
  wire [26:0] n421_o;
  wire n423_o;
  wire [26:0] n424_o;
  reg [26:0] n425_o;
  wire [24:0] n426_o;
  wire [26:0] n428_o;
  wire [5:0] n429_o;
  wire [2:0] n430_o;
  wire [8:0] n431_o;
  wire [2:0] selfunctiontable10_n432;
  wire [2:0] selfunctiontable10_y;
  wire [26:0] n436_o;
  wire n438_o;
  wire n440_o;
  wire n441_o;
  wire [25:0] n443_o;
  wire [26:0] n445_o;
  wire n447_o;
  wire n449_o;
  wire n450_o;
  wire [1:0] n452_o;
  reg [26:0] n453_o;
  wire n454_o;
  wire [26:0] n455_o;
  wire n457_o;
  wire [26:0] n458_o;
  reg [26:0] n459_o;
  wire [24:0] n460_o;
  wire [26:0] n462_o;
  wire [5:0] n463_o;
  wire [2:0] n464_o;
  wire [8:0] n465_o;
  wire [2:0] selfunctiontable9_n466;
  wire [2:0] selfunctiontable9_y;
  wire [26:0] n470_o;
  wire n472_o;
  wire n474_o;
  wire n475_o;
  wire [25:0] n477_o;
  wire [26:0] n479_o;
  wire n481_o;
  wire n483_o;
  wire n484_o;
  wire [1:0] n486_o;
  reg [26:0] n487_o;
  wire n488_o;
  wire [26:0] n489_o;
  wire n491_o;
  wire [26:0] n492_o;
  reg [26:0] n493_o;
  wire [24:0] n494_o;
  wire [26:0] n496_o;
  wire [5:0] n497_o;
  wire [2:0] n498_o;
  wire [8:0] n499_o;
  wire [2:0] selfunctiontable8_n500;
  wire [2:0] selfunctiontable8_y;
  wire [26:0] n504_o;
  wire n506_o;
  wire n508_o;
  wire n509_o;
  wire [25:0] n511_o;
  wire [26:0] n513_o;
  wire n515_o;
  wire n517_o;
  wire n518_o;
  wire [1:0] n520_o;
  reg [26:0] n521_o;
  wire n522_o;
  wire [26:0] n523_o;
  wire n525_o;
  wire [26:0] n526_o;
  reg [26:0] n527_o;
  wire [24:0] n528_o;
  wire [26:0] n530_o;
  wire [5:0] n531_o;
  wire [2:0] n532_o;
  wire [8:0] n533_o;
  wire [2:0] selfunctiontable7_n534;
  wire [2:0] selfunctiontable7_y;
  wire [26:0] n538_o;
  wire n540_o;
  wire n542_o;
  wire n543_o;
  wire [25:0] n545_o;
  wire [26:0] n547_o;
  wire n549_o;
  wire n551_o;
  wire n552_o;
  wire [1:0] n554_o;
  reg [26:0] n555_o;
  wire n556_o;
  wire [26:0] n557_o;
  wire n559_o;
  wire [26:0] n560_o;
  reg [26:0] n561_o;
  wire [24:0] n562_o;
  wire [26:0] n564_o;
  wire [5:0] n565_o;
  wire [2:0] n566_o;
  wire [8:0] n567_o;
  wire [2:0] selfunctiontable6_n568;
  wire [2:0] selfunctiontable6_y;
  wire [26:0] n572_o;
  wire n574_o;
  wire n576_o;
  wire n577_o;
  wire [25:0] n579_o;
  wire [26:0] n581_o;
  wire n583_o;
  wire n585_o;
  wire n586_o;
  wire [1:0] n588_o;
  reg [26:0] n589_o;
  wire n590_o;
  wire [26:0] n591_o;
  wire n593_o;
  wire [26:0] n594_o;
  reg [26:0] n595_o;
  wire [24:0] n596_o;
  wire [26:0] n598_o;
  wire [5:0] n599_o;
  wire [2:0] n600_o;
  wire [8:0] n601_o;
  wire [2:0] selfunctiontable5_n602;
  wire [2:0] selfunctiontable5_y;
  wire [26:0] n606_o;
  wire n608_o;
  wire n610_o;
  wire n611_o;
  wire [25:0] n613_o;
  wire [26:0] n615_o;
  wire n617_o;
  wire n619_o;
  wire n620_o;
  wire [1:0] n622_o;
  reg [26:0] n623_o;
  wire n624_o;
  wire [26:0] n625_o;
  wire n627_o;
  wire [26:0] n628_o;
  reg [26:0] n629_o;
  wire [24:0] n630_o;
  wire [26:0] n632_o;
  wire [5:0] n633_o;
  wire [2:0] n634_o;
  wire [8:0] n635_o;
  wire [2:0] selfunctiontable4_n636;
  wire [2:0] selfunctiontable4_y;
  wire [26:0] n640_o;
  wire n642_o;
  wire n644_o;
  wire n645_o;
  wire [25:0] n647_o;
  wire [26:0] n649_o;
  wire n651_o;
  wire n653_o;
  wire n654_o;
  wire [1:0] n656_o;
  reg [26:0] n657_o;
  wire n658_o;
  wire [26:0] n659_o;
  wire n661_o;
  wire [26:0] n662_o;
  reg [26:0] n663_o;
  wire [24:0] n664_o;
  wire [26:0] n666_o;
  wire [5:0] n667_o;
  wire [2:0] n668_o;
  wire [8:0] n669_o;
  wire [2:0] selfunctiontable3_n670;
  wire [2:0] selfunctiontable3_y;
  wire [26:0] n674_o;
  wire n676_o;
  wire n678_o;
  wire n679_o;
  wire [25:0] n681_o;
  wire [26:0] n683_o;
  wire n685_o;
  wire n687_o;
  wire n688_o;
  wire [1:0] n690_o;
  reg [26:0] n691_o;
  wire n692_o;
  wire [26:0] n693_o;
  wire n695_o;
  wire [26:0] n696_o;
  reg [26:0] n697_o;
  wire [24:0] n698_o;
  wire [26:0] n700_o;
  wire [5:0] n701_o;
  wire [2:0] n702_o;
  wire [8:0] n703_o;
  wire [2:0] selfunctiontable2_n704;
  wire [2:0] selfunctiontable2_y;
  wire [26:0] n708_o;
  wire n710_o;
  wire n712_o;
  wire n713_o;
  wire [25:0] n715_o;
  wire [26:0] n717_o;
  wire n719_o;
  wire n721_o;
  wire n722_o;
  wire [1:0] n724_o;
  reg [26:0] n725_o;
  wire n726_o;
  wire [26:0] n727_o;
  wire n729_o;
  wire [26:0] n730_o;
  reg [26:0] n731_o;
  wire [24:0] n732_o;
  wire [26:0] n734_o;
  wire [5:0] n735_o;
  wire [2:0] n736_o;
  wire [8:0] n737_o;
  wire [2:0] selfunctiontable1_n738;
  wire [2:0] selfunctiontable1_y;
  wire [26:0] n742_o;
  wire n744_o;
  wire n746_o;
  wire n747_o;
  wire [25:0] n749_o;
  wire [26:0] n751_o;
  wire n753_o;
  wire n755_o;
  wire n756_o;
  wire [1:0] n758_o;
  reg [26:0] n759_o;
  wire n760_o;
  wire [26:0] n761_o;
  wire n763_o;
  wire [26:0] n764_o;
  reg [26:0] n765_o;
  wire [24:0] n766_o;
  wire n767_o;
  wire [1:0] n768_o;
  wire n769_o;
  wire [1:0] n771_o;
  wire [1:0] n772_o;
  wire n773_o;
  wire [1:0] n775_o;
  wire [1:0] n776_o;
  wire n777_o;
  wire [1:0] n779_o;
  wire [1:0] n780_o;
  wire n781_o;
  wire [1:0] n783_o;
  wire [1:0] n784_o;
  wire n785_o;
  wire [1:0] n787_o;
  wire [1:0] n788_o;
  wire n789_o;
  wire [1:0] n791_o;
  wire [1:0] n792_o;
  wire n793_o;
  wire [1:0] n795_o;
  wire [1:0] n796_o;
  wire n797_o;
  wire [1:0] n799_o;
  wire [1:0] n800_o;
  wire n801_o;
  wire [1:0] n803_o;
  wire [1:0] n804_o;
  wire n805_o;
  wire [1:0] n807_o;
  wire [1:0] n808_o;
  wire n809_o;
  wire [1:0] n811_o;
  wire [1:0] n812_o;
  wire n813_o;
  wire [1:0] n815_o;
  wire [1:0] n816_o;
  wire n817_o;
  wire [1:0] n819_o;
  wire [1:0] n820_o;
  wire n821_o;
  wire [1:0] n823_o;
  wire [3:0] n824_o;
  wire [5:0] n825_o;
  wire [7:0] n826_o;
  wire [9:0] n827_o;
  wire [11:0] n828_o;
  wire [13:0] n829_o;
  wire [15:0] n830_o;
  wire [17:0] n831_o;
  wire [19:0] n832_o;
  wire [21:0] n833_o;
  wire [23:0] n834_o;
  wire [25:0] n835_o;
  wire [27:0] n836_o;
  wire n837_o;
  wire [2:0] n838_o;
  wire [4:0] n839_o;
  wire [6:0] n840_o;
  wire [8:0] n841_o;
  wire [10:0] n842_o;
  wire [12:0] n843_o;
  wire [14:0] n844_o;
  wire [16:0] n845_o;
  wire [18:0] n846_o;
  wire [20:0] n847_o;
  wire [22:0] n848_o;
  wire [24:0] n849_o;
  wire [26:0] n850_o;
  wire [27:0] n851_o;
  wire [27:0] n852_o;
  wire [25:0] n853_o;
  wire [23:0] n854_o;
  wire n855_o;
  wire [23:0] n856_o;
  wire [23:0] n857_o;
  wire n858_o;
  wire n859_o;
  wire [9:0] n861_o;
  wire [9:0] n862_o;
  wire [22:0] n863_o;
  wire [32:0] n864_o;
  wire [32:0] n866_o;
  wire [32:0] n867_o;
  wire n869_o;
  wire [1:0] n870_o;
  wire [1:0] n872_o;
  wire n874_o;
  wire [1:0] n875_o;
  wire n878_o;
  reg [1:0] n879_o;
  wire [2:0] n880_o;
  wire [30:0] n881_o;
  wire [33:0] n882_o;
  reg [9:0] n883_q;
  reg [9:0] n884_q;
  reg [9:0] n885_q;
  reg [9:0] n886_q;
  reg [9:0] n887_q;
  reg [9:0] n888_q;
  reg [9:0] n889_q;
  reg [9:0] n890_q;
  reg [9:0] n891_q;
  reg [9:0] n892_q;
  reg [9:0] n893_q;
  reg [9:0] n894_q;
  reg n895_q;
  reg n896_q;
  reg n897_q;
  reg n898_q;
  reg n899_q;
  reg n900_q;
  reg n901_q;
  reg n902_q;
  reg n903_q;
  reg n904_q;
  reg n905_q;
  reg n906_q;
  reg [1:0] n907_q;
  reg [1:0] n908_q;
  reg [1:0] n909_q;
  reg [1:0] n910_q;
  reg [1:0] n911_q;
  reg [1:0] n912_q;
  reg [1:0] n913_q;
  reg [1:0] n914_q;
  reg [1:0] n915_q;
  reg [1:0] n916_q;
  reg [1:0] n917_q;
  reg [1:0] n918_q;
  reg [23:0] n919_q;
  reg [23:0] n920_q;
  reg [23:0] n921_q;
  reg [23:0] n922_q;
  reg [23:0] n923_q;
  reg [23:0] n924_q;
  reg [23:0] n925_q;
  reg [23:0] n926_q;
  reg [23:0] n927_q;
  reg [23:0] n928_q;
  reg [23:0] n929_q;
  reg [26:0] n930_q;
  reg [2:0] n931_q;
  reg [26:0] n932_q;
  reg [2:0] n933_q;
  reg [26:0] n934_q;
  reg [2:0] n935_q;
  reg [26:0] n936_q;
  reg [2:0] n937_q;
  reg [26:0] n938_q;
  reg [26:0] n939_q;
  reg [2:0] n940_q;
  reg [26:0] n941_q;
  reg [26:0] n942_q;
  reg [2:0] n943_q;
  reg [26:0] n944_q;
  reg [26:0] n945_q;
  reg [2:0] n946_q;
  reg [26:0] n947_q;
  reg [2:0] n948_q;
  reg [26:0] n949_q;
  reg [2:0] n950_q;
  reg [26:0] n951_q;
  reg [2:0] n952_q;
  reg [26:0] n953_q;
  reg [2:0] n954_q;
  reg [26:0] n955_q;
  reg [26:0] n956_q;
  reg [2:0] n957_q;
  reg [26:0] n958_q;
  reg [1:0] n959_q;
  reg [1:0] n960_q;
  reg [1:0] n961_q;
  reg [1:0] n962_q;
  reg [1:0] n963_q;
  reg [1:0] n964_q;
  reg [1:0] n965_q;
  reg [1:0] n966_q;
  reg [1:0] n967_q;
  reg [1:0] n968_q;
  reg [1:0] n969_q;
  reg [1:0] n970_q;
  reg [1:0] n971_q;
  reg [1:0] n972_q;
  reg [1:0] n973_q;
  reg [1:0] n974_q;
  reg [1:0] n975_q;
  reg [1:0] n976_q;
  reg [1:0] n977_q;
  reg [1:0] n978_q;
  reg [1:0] n979_q;
  reg [1:0] n980_q;
  reg [1:0] n981_q;
  reg [1:0] n982_q;
  reg [1:0] n983_q;
  reg [1:0] n984_q;
  reg [1:0] n985_q;
  reg [1:0] n986_q;
  reg [1:0] n987_q;
  reg [1:0] n988_q;
  reg [1:0] n989_q;
  reg [1:0] n990_q;
  reg [1:0] n991_q;
  reg [1:0] n992_q;
  reg [1:0] n993_q;
  reg [1:0] n994_q;
  reg [1:0] n995_q;
  reg [1:0] n996_q;
  reg [1:0] n997_q;
  reg [1:0] n998_q;
  reg [1:0] n999_q;
  reg [1:0] n1000_q;
  reg [1:0] n1001_q;
  reg [1:0] n1002_q;
  reg [1:0] n1003_q;
  reg [1:0] n1004_q;
  reg [1:0] n1005_q;
  reg [1:0] n1006_q;
  reg [1:0] n1007_q;
  reg [1:0] n1008_q;
  reg [1:0] n1009_q;
  reg [1:0] n1010_q;
  reg [1:0] n1011_q;
  reg [1:0] n1012_q;
  reg [1:0] n1013_q;
  reg [1:0] n1014_q;
  reg [1:0] n1015_q;
  reg [1:0] n1016_q;
  reg [1:0] n1017_q;
  reg [1:0] n1018_q;
  reg [1:0] n1019_q;
  reg [1:0] n1020_q;
  reg [1:0] n1021_q;
  reg [1:0] n1022_q;
  reg [1:0] n1023_q;
  reg [1:0] n1024_q;
  reg [1:0] n1025_q;
  reg [1:0] n1026_q;
  reg [1:0] n1027_q;
  reg [1:0] n1028_q;
  reg [1:0] n1029_q;
  reg [1:0] n1030_q;
  reg [1:0] n1031_q;
  reg [1:0] n1032_q;
  reg [1:0] n1033_q;
  reg [1:0] n1034_q;
  reg [1:0] n1035_q;
  reg [1:0] n1036_q;
  reg [1:0] n1037_q;
  reg [1:0] n1038_q;
  reg [1:0] n1039_q;
  reg [1:0] n1040_q;
  reg [1:0] n1041_q;
  reg [1:0] n1042_q;
  reg [1:0] n1043_q;
  reg [1:0] n1044_q;
  reg [1:0] n1045_q;
  reg [1:0] n1046_q;
  reg [1:0] n1047_q;
  reg [1:0] n1048_q;
  reg [1:0] n1049_q;
  reg [1:0] n1050_q;
  reg [1:0] n1051_q;
  reg [1:0] n1052_q;
  reg [1:0] n1053_q;
  reg [1:0] n1054_q;
  reg [1:0] n1055_q;
  reg [1:0] n1056_q;
  reg [1:0] n1057_q;
  reg [1:0] n1058_q;
  reg [1:0] n1059_q;
  reg [1:0] n1060_q;
  reg [1:0] n1061_q;
  reg [1:0] n1062_q;
  reg [1:0] n1063_q;
  reg [1:0] n1064_q;
  reg [1:0] n1065_q;
  reg [1:0] n1066_q;
  reg [1:0] n1067_q;
  reg [1:0] n1068_q;
  reg [1:0] n1069_q;
  reg [1:0] n1070_q;
  reg [1:0] n1071_q;
  reg [1:0] n1072_q;
  reg [1:0] n1073_q;
  reg [1:0] n1074_q;
  reg [1:0] n1075_q;
  reg [1:0] n1076_q;
  reg [1:0] n1077_q;
  reg [1:0] n1078_q;
  reg [1:0] n1079_q;
  reg [1:0] n1080_q;
  reg [1:0] n1081_q;
  reg [1:0] n1082_q;
  reg [1:0] n1083_q;
  reg [1:0] n1084_q;
  reg [1:0] n1085_q;
  reg [1:0] n1086_q;
  reg [1:0] n1087_q;
  reg [1:0] n1088_q;
  reg [1:0] n1089_q;
  reg [1:0] n1090_q;
  reg [1:0] n1091_q;
  reg [1:0] n1092_q;
  reg [1:0] n1093_q;
  reg [1:0] n1094_q;
  reg [1:0] n1095_q;
  reg [1:0] n1096_q;
  reg [1:0] n1097_q;
  reg [1:0] n1098_q;
  reg [1:0] n1099_q;
  reg [1:0] n1100_q;
  reg [1:0] n1101_q;
  reg [1:0] n1102_q;
  reg [1:0] n1103_q;
  reg [1:0] n1104_q;
  reg [1:0] n1105_q;
  reg [1:0] n1106_q;
  reg [1:0] n1107_q;
  reg [1:0] n1108_q;
  reg [1:0] n1109_q;
  reg [1:0] n1110_q;
  reg [1:0] n1111_q;
  reg [1:0] n1112_q;
  reg [1:0] n1113_q;
  reg [1:0] n1114_q;
  reg [1:0] n1115_q;
  reg [1:0] n1116_q;
  reg [1:0] n1117_q;
  reg [1:0] n1118_q;
  reg [1:0] n1119_q;
  reg [1:0] n1120_q;
  reg [1:0] n1121_q;
  reg [1:0] n1122_q;
  reg [27:0] n1123_q;
  assign R = n882_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:588:8  */
  assign fx = n248_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:589:8  */
  assign fy = n251_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:8  */
  assign expr0 = n258_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:15  */
  assign expr0_d1 = n883_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:25  */
  assign expr0_d2 = n884_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:35  */
  assign expr0_d3 = n885_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:45  */
  assign expr0_d4 = n886_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:55  */
  assign expr0_d5 = n887_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:65  */
  assign expr0_d6 = n888_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:75  */
  assign expr0_d7 = n889_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:85  */
  assign expr0_d8 = n890_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:95  */
  assign expr0_d9 = n891_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:105  */
  assign expr0_d10 = n892_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:116  */
  assign expr0_d11 = n893_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:590:127  */
  assign expr0_d12 = n894_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:8  */
  assign sr = n261_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:12  */
  assign sr_d1 = n895_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:19  */
  assign sr_d2 = n896_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:26  */
  assign sr_d3 = n897_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:33  */
  assign sr_d4 = n898_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:40  */
  assign sr_d5 = n899_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:47  */
  assign sr_d6 = n900_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:54  */
  assign sr_d7 = n901_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:61  */
  assign sr_d8 = n902_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:68  */
  assign sr_d9 = n903_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:75  */
  assign sr_d10 = n904_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:83  */
  assign sr_d11 = n905_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:591:91  */
  assign sr_d12 = n906_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:592:8  */
  assign exnxy = n264_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:8  */
  assign exnr0 = n288_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:15  */
  assign exnr0_d1 = n907_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:25  */
  assign exnr0_d2 = n908_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:35  */
  assign exnr0_d3 = n909_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:45  */
  assign exnr0_d4 = n910_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:55  */
  assign exnr0_d5 = n911_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:65  */
  assign exnr0_d6 = n912_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:75  */
  assign exnr0_d7 = n913_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:85  */
  assign exnr0_d8 = n914_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:95  */
  assign exnr0_d9 = n915_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:105  */
  assign exnr0_d10 = n916_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:116  */
  assign exnr0_d11 = n917_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:593:127  */
  assign exnr0_d12 = n918_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:8  */
  assign d = fy; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:11  */
  assign d_d1 = n919_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:17  */
  assign d_d2 = n920_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:23  */
  assign d_d3 = n921_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:29  */
  assign d_d4 = n922_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:35  */
  assign d_d5 = n923_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:41  */
  assign d_d6 = n924_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:47  */
  assign d_d7 = n925_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:53  */
  assign d_d8 = n926_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:59  */
  assign d_d9 = n927_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:65  */
  assign d_d10 = n928_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:594:72  */
  assign d_d11 = n929_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:595:8  */
  assign psx = n290_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:596:8  */
  assign betaw14 = n292_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:597:8  */
  assign sel14 = n295_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:598:8  */
  assign q14 = q14_copy5; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:599:8  */
  assign q14_copy5 = selfunctiontable14_n296; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:600:8  */
  assign absq14d = n317_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:601:8  */
  assign w13 = n323_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:602:8  */
  assign betaw13 = n326_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:602:17  */
  assign betaw13_d1 = n930_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:603:8  */
  assign sel13 = n329_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:604:8  */
  assign q13 = q13_copy6_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:605:8  */
  assign q13_copy6 = selfunctiontable13_n330; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:605:19  */
  assign q13_copy6_d1 = n931_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:606:8  */
  assign absq13d = n351_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:607:8  */
  assign w12 = n357_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:608:8  */
  assign betaw12 = n360_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:608:17  */
  assign betaw12_d1 = n932_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:609:8  */
  assign sel12 = n363_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:610:8  */
  assign q12 = q12_copy7_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:611:8  */
  assign q12_copy7 = selfunctiontable12_n364; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:611:19  */
  assign q12_copy7_d1 = n933_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:612:8  */
  assign absq12d = n385_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:613:8  */
  assign w11 = n391_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:614:8  */
  assign betaw11 = n394_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:614:17  */
  assign betaw11_d1 = n934_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:615:8  */
  assign sel11 = n397_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:616:8  */
  assign q11 = q11_copy8_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:617:8  */
  assign q11_copy8 = selfunctiontable11_n398; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:617:19  */
  assign q11_copy8_d1 = n935_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:618:8  */
  assign absq11d = n419_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:619:8  */
  assign w10 = n425_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:620:8  */
  assign betaw10 = n428_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:620:17  */
  assign betaw10_d1 = n936_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:621:8  */
  assign sel10 = n431_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:622:8  */
  assign q10 = q10_copy9; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:622:13  */
  assign q10_d1 = n937_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:623:8  */
  assign q10_copy9 = selfunctiontable10_n432; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:624:8  */
  assign absq10d = n453_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:624:17  */
  assign absq10d_d1 = n938_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:625:8  */
  assign w9 = n459_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:626:8  */
  assign betaw9 = n462_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:626:16  */
  assign betaw9_d1 = n939_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:627:8  */
  assign sel9 = n465_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:628:8  */
  assign q9 = q9_copy10; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:628:12  */
  assign q9_d1 = n940_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:629:8  */
  assign q9_copy10 = selfunctiontable9_n466; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:630:8  */
  assign absq9d = n487_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:630:16  */
  assign absq9d_d1 = n941_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:631:8  */
  assign w8 = n493_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:632:8  */
  assign betaw8 = n496_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:632:16  */
  assign betaw8_d1 = n942_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:633:8  */
  assign sel8 = n499_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:634:8  */
  assign q8 = q8_copy11; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:634:12  */
  assign q8_d1 = n943_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:635:8  */
  assign q8_copy11 = selfunctiontable8_n500; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:636:8  */
  assign absq8d = n521_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:636:16  */
  assign absq8d_d1 = n944_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:637:8  */
  assign w7 = n527_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:638:8  */
  assign betaw7 = n530_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:639:8  */
  assign sel7 = n533_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:640:8  */
  assign q7 = q7_copy12; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:641:8  */
  assign q7_copy12 = selfunctiontable7_n534; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:642:8  */
  assign absq7d = n555_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:643:8  */
  assign w6 = n561_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:644:8  */
  assign betaw6 = n564_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:644:16  */
  assign betaw6_d1 = n945_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:645:8  */
  assign sel6 = n567_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:646:8  */
  assign q6 = q6_copy13_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:647:8  */
  assign q6_copy13 = selfunctiontable6_n568; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:647:19  */
  assign q6_copy13_d1 = n946_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:648:8  */
  assign absq6d = n589_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:649:8  */
  assign w5 = n595_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:650:8  */
  assign betaw5 = n598_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:650:16  */
  assign betaw5_d1 = n947_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:651:8  */
  assign sel5 = n601_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:652:8  */
  assign q5 = q5_copy14_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:653:8  */
  assign q5_copy14 = selfunctiontable5_n602; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:653:19  */
  assign q5_copy14_d1 = n948_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:654:8  */
  assign absq5d = n623_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:655:8  */
  assign w4 = n629_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:656:8  */
  assign betaw4 = n632_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:656:16  */
  assign betaw4_d1 = n949_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:657:8  */
  assign sel4 = n635_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:658:8  */
  assign q4 = q4_copy15_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:659:8  */
  assign q4_copy15 = selfunctiontable4_n636; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:659:19  */
  assign q4_copy15_d1 = n950_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:660:8  */
  assign absq4d = n657_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:661:8  */
  assign w3 = n663_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:662:8  */
  assign betaw3 = n666_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:662:16  */
  assign betaw3_d1 = n951_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:663:8  */
  assign sel3 = n669_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:664:8  */
  assign q3 = q3_copy16_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:665:8  */
  assign q3_copy16 = selfunctiontable3_n670; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:665:19  */
  assign q3_copy16_d1 = n952_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:666:8  */
  assign absq3d = n691_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:667:8  */
  assign w2 = n697_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:668:8  */
  assign betaw2 = n700_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:668:16  */
  assign betaw2_d1 = n953_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:669:8  */
  assign sel2 = n703_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:670:8  */
  assign q2 = q2_copy17; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:670:12  */
  assign q2_d1 = n954_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:671:8  */
  assign q2_copy17 = selfunctiontable2_n704; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:672:8  */
  assign absq2d = n725_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:672:16  */
  assign absq2d_d1 = n955_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:673:8  */
  assign w1 = n731_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:674:8  */
  assign betaw1 = n734_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:674:16  */
  assign betaw1_d1 = n956_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:675:8  */
  assign sel1 = n737_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:676:8  */
  assign q1 = q1_copy18; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:676:12  */
  assign q1_d1 = n957_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:677:8  */
  assign q1_copy18 = selfunctiontable1_n738; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:678:8  */
  assign absq1d = n759_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:678:16  */
  assign absq1d_d1 = n958_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:679:8  */
  assign w0 = n765_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:680:8  */
  assign wfinal = n766_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:681:8  */
  assign qm0 = n767_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:8  */
  assign qp14 = n768_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:14  */
  assign qp14_d1 = n959_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:23  */
  assign qp14_d2 = n960_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:32  */
  assign qp14_d3 = n961_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:41  */
  assign qp14_d4 = n962_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:50  */
  assign qp14_d5 = n963_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:59  */
  assign qp14_d6 = n964_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:68  */
  assign qp14_d7 = n965_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:77  */
  assign qp14_d8 = n966_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:86  */
  assign qp14_d9 = n967_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:95  */
  assign qp14_d10 = n968_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:682:105  */
  assign qp14_d11 = n969_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:8  */
  assign qm14 = n771_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:14  */
  assign qm14_d1 = n970_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:23  */
  assign qm14_d2 = n971_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:32  */
  assign qm14_d3 = n972_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:41  */
  assign qm14_d4 = n973_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:50  */
  assign qm14_d5 = n974_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:59  */
  assign qm14_d6 = n975_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:68  */
  assign qm14_d7 = n976_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:77  */
  assign qm14_d8 = n977_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:86  */
  assign qm14_d9 = n978_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:95  */
  assign qm14_d10 = n979_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:105  */
  assign qm14_d11 = n980_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:683:115  */
  assign qm14_d12 = n981_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:8  */
  assign qp13 = n772_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:14  */
  assign qp13_d1 = n982_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:23  */
  assign qp13_d2 = n983_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:32  */
  assign qp13_d3 = n984_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:41  */
  assign qp13_d4 = n985_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:50  */
  assign qp13_d5 = n986_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:59  */
  assign qp13_d6 = n987_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:68  */
  assign qp13_d7 = n988_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:77  */
  assign qp13_d8 = n989_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:86  */
  assign qp13_d9 = n990_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:684:95  */
  assign qp13_d10 = n991_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:8  */
  assign qm13 = n775_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:14  */
  assign qm13_d1 = n992_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:23  */
  assign qm13_d2 = n993_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:32  */
  assign qm13_d3 = n994_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:41  */
  assign qm13_d4 = n995_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:50  */
  assign qm13_d5 = n996_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:59  */
  assign qm13_d6 = n997_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:68  */
  assign qm13_d7 = n998_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:77  */
  assign qm13_d8 = n999_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:86  */
  assign qm13_d9 = n1000_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:95  */
  assign qm13_d10 = n1001_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:685:105  */
  assign qm13_d11 = n1002_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:8  */
  assign qp12 = n776_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:14  */
  assign qp12_d1 = n1003_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:23  */
  assign qp12_d2 = n1004_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:32  */
  assign qp12_d3 = n1005_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:41  */
  assign qp12_d4 = n1006_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:50  */
  assign qp12_d5 = n1007_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:59  */
  assign qp12_d6 = n1008_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:68  */
  assign qp12_d7 = n1009_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:77  */
  assign qp12_d8 = n1010_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:686:86  */
  assign qp12_d9 = n1011_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:8  */
  assign qm12 = n779_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:14  */
  assign qm12_d1 = n1012_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:23  */
  assign qm12_d2 = n1013_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:32  */
  assign qm12_d3 = n1014_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:41  */
  assign qm12_d4 = n1015_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:50  */
  assign qm12_d5 = n1016_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:59  */
  assign qm12_d6 = n1017_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:68  */
  assign qm12_d7 = n1018_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:77  */
  assign qm12_d8 = n1019_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:86  */
  assign qm12_d9 = n1020_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:687:95  */
  assign qm12_d10 = n1021_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:8  */
  assign qp11 = n780_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:14  */
  assign qp11_d1 = n1022_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:23  */
  assign qp11_d2 = n1023_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:32  */
  assign qp11_d3 = n1024_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:41  */
  assign qp11_d4 = n1025_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:50  */
  assign qp11_d5 = n1026_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:59  */
  assign qp11_d6 = n1027_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:68  */
  assign qp11_d7 = n1028_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:688:77  */
  assign qp11_d8 = n1029_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:8  */
  assign qm11 = n783_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:14  */
  assign qm11_d1 = n1030_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:23  */
  assign qm11_d2 = n1031_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:32  */
  assign qm11_d3 = n1032_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:41  */
  assign qm11_d4 = n1033_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:50  */
  assign qm11_d5 = n1034_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:59  */
  assign qm11_d6 = n1035_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:68  */
  assign qm11_d7 = n1036_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:77  */
  assign qm11_d8 = n1037_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:689:86  */
  assign qm11_d9 = n1038_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:8  */
  assign qp10 = n784_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:14  */
  assign qp10_d1 = n1039_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:23  */
  assign qp10_d2 = n1040_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:32  */
  assign qp10_d3 = n1041_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:41  */
  assign qp10_d4 = n1042_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:50  */
  assign qp10_d5 = n1043_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:59  */
  assign qp10_d6 = n1044_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:68  */
  assign qp10_d7 = n1045_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:690:77  */
  assign qp10_d8 = n1046_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:8  */
  assign qm10 = n787_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:14  */
  assign qm10_d1 = n1047_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:23  */
  assign qm10_d2 = n1048_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:32  */
  assign qm10_d3 = n1049_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:41  */
  assign qm10_d4 = n1050_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:50  */
  assign qm10_d5 = n1051_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:59  */
  assign qm10_d6 = n1052_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:68  */
  assign qm10_d7 = n1053_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:77  */
  assign qm10_d8 = n1054_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:691:86  */
  assign qm10_d9 = n1055_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:8  */
  assign qp9 = n788_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:13  */
  assign qp9_d1 = n1056_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:21  */
  assign qp9_d2 = n1057_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:29  */
  assign qp9_d3 = n1058_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:37  */
  assign qp9_d4 = n1059_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:45  */
  assign qp9_d5 = n1060_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:53  */
  assign qp9_d6 = n1061_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:692:61  */
  assign qp9_d7 = n1062_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:8  */
  assign qm9 = n791_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:13  */
  assign qm9_d1 = n1063_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:21  */
  assign qm9_d2 = n1064_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:29  */
  assign qm9_d3 = n1065_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:37  */
  assign qm9_d4 = n1066_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:45  */
  assign qm9_d5 = n1067_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:53  */
  assign qm9_d6 = n1068_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:61  */
  assign qm9_d7 = n1069_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:693:69  */
  assign qm9_d8 = n1070_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:8  */
  assign qp8 = n792_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:13  */
  assign qp8_d1 = n1071_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:21  */
  assign qp8_d2 = n1072_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:29  */
  assign qp8_d3 = n1073_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:37  */
  assign qp8_d4 = n1074_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:45  */
  assign qp8_d5 = n1075_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:694:53  */
  assign qp8_d6 = n1076_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:8  */
  assign qm8 = n795_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:13  */
  assign qm8_d1 = n1077_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:21  */
  assign qm8_d2 = n1078_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:29  */
  assign qm8_d3 = n1079_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:37  */
  assign qm8_d4 = n1080_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:45  */
  assign qm8_d5 = n1081_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:53  */
  assign qm8_d6 = n1082_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:695:61  */
  assign qm8_d7 = n1083_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:8  */
  assign qp7 = n796_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:13  */
  assign qp7_d1 = n1084_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:21  */
  assign qp7_d2 = n1085_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:29  */
  assign qp7_d3 = n1086_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:37  */
  assign qp7_d4 = n1087_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:696:45  */
  assign qp7_d5 = n1088_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:8  */
  assign qm7 = n799_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:13  */
  assign qm7_d1 = n1089_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:21  */
  assign qm7_d2 = n1090_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:29  */
  assign qm7_d3 = n1091_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:37  */
  assign qm7_d4 = n1092_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:45  */
  assign qm7_d5 = n1093_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:697:53  */
  assign qm7_d6 = n1094_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:698:8  */
  assign qp6 = n800_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:698:13  */
  assign qp6_d1 = n1095_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:698:21  */
  assign qp6_d2 = n1096_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:698:29  */
  assign qp6_d3 = n1097_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:698:37  */
  assign qp6_d4 = n1098_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:8  */
  assign qm6 = n803_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:13  */
  assign qm6_d1 = n1099_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:21  */
  assign qm6_d2 = n1100_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:29  */
  assign qm6_d3 = n1101_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:37  */
  assign qm6_d4 = n1102_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:699:45  */
  assign qm6_d5 = n1103_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:700:8  */
  assign qp5 = n804_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:700:13  */
  assign qp5_d1 = n1104_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:700:21  */
  assign qp5_d2 = n1105_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:700:29  */
  assign qp5_d3 = n1106_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:701:8  */
  assign qm5 = n807_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:701:13  */
  assign qm5_d1 = n1107_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:701:21  */
  assign qm5_d2 = n1108_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:701:29  */
  assign qm5_d3 = n1109_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:701:37  */
  assign qm5_d4 = n1110_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:702:8  */
  assign qp4 = n808_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:702:13  */
  assign qp4_d1 = n1111_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:702:21  */
  assign qp4_d2 = n1112_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:703:8  */
  assign qm4 = n811_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:703:13  */
  assign qm4_d1 = n1113_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:703:21  */
  assign qm4_d2 = n1114_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:703:29  */
  assign qm4_d3 = n1115_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:704:8  */
  assign qp3 = n812_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:704:13  */
  assign qp3_d1 = n1116_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:705:8  */
  assign qm3 = n815_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:705:13  */
  assign qm3_d1 = n1117_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:705:21  */
  assign qm3_d2 = n1118_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:706:8  */
  assign qp2 = n816_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:706:13  */
  assign qp2_d1 = n1119_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:707:8  */
  assign qm2 = n819_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:707:13  */
  assign qm2_d1 = n1120_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:707:21  */
  assign qm2_d2 = n1121_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:708:8  */
  assign qp1 = n820_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:709:8  */
  assign qm1 = n823_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:709:13  */
  assign qm1_d1 = n1122_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:710:8  */
  assign qp = n836_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:710:12  */
  assign qp_d1 = n1123_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:711:8  */
  assign qm = n851_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:712:8  */
  assign quotient = n852_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:713:8  */
  assign mr = n853_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:714:8  */
  assign frnorm = n856_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:715:8  */
  assign round = n858_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:716:8  */
  assign expr1 = n862_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:717:8  */
  assign expfrac = n864_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:718:8  */
  assign expfracr = n867_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:719:8  */
  assign exnr = n870_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:720:8  */
  assign exnrfinal = n879_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:968:17  */
  assign n246_o = X[22:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:968:14  */
  assign n248_o = {1'b1, n246_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:969:17  */
  assign n249_o = Y[22:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:969:14  */
  assign n251_o = {1'b1, n249_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:971:22  */
  assign n252_o = X[30:23];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:971:19  */
  assign n254_o = {2'b00, n252_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:971:49  */
  assign n255_o = Y[30:23];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:971:46  */
  assign n257_o = {2'b00, n255_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:971:38  */
  assign n258_o = n254_o - n257_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:972:11  */
  assign n259_o = X[31];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:972:21  */
  assign n260_o = Y[31];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:972:16  */
  assign n261_o = n259_o ^ n260_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:974:14  */
  assign n262_o = X[33:32];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:974:32  */
  assign n263_o = Y[33:32];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:974:29  */
  assign n264_o = {n262_o, n263_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:977:18  */
  assign n267_o = exnxy == 4'b0101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:978:18  */
  assign n270_o = exnxy == 4'b0001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:978:30  */
  assign n272_o = exnxy == 4'b0010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:978:30  */
  assign n273_o = n270_o | n272_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:978:39  */
  assign n275_o = exnxy == 4'b0110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:978:39  */
  assign n276_o = n273_o | n275_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:979:18  */
  assign n279_o = exnxy == 4'b0100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:979:30  */
  assign n281_o = exnxy == 4'b1000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:979:30  */
  assign n282_o = n279_o | n281_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:979:39  */
  assign n284_o = exnxy == 4'b1001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:979:39  */
  assign n285_o = n282_o | n284_o;
  assign n287_o = {n285_o, n276_o, n267_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:975:4  */
  always @*
    case (n287_o)
      3'b100: n288_o = 2'b10;
      3'b010: n288_o = 2'b00;
      3'b001: n288_o = 2'b01;
      default: n288_o = 2'b11;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:982:15  */
  assign n290_o = {1'b0, fx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:983:21  */
  assign n292_o = {2'b00, psx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:984:20  */
  assign n293_o = betaw14[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:984:38  */
  assign n294_o = d[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:984:35  */
  assign n295_o = {n293_o, n294_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:987:23  */
  assign selfunctiontable14_n296 = selfunctiontable14_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:985:4  */
  selfunction_f300_uid4 selfunctiontable14 (
    .x(sel14),
    .y(selfunctiontable14_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:992:16  */
  assign n300_o = {3'b000, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:992:66  */
  assign n302_o = q14 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:992:77  */
  assign n304_o = q14 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:992:77  */
  assign n305_o = n302_o | n304_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:993:15  */
  assign n307_o = {2'b00, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:993:19  */
  assign n309_o = {n307_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:993:52  */
  assign n311_o = q14 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:993:63  */
  assign n313_o = q14 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:993:63  */
  assign n314_o = n311_o | n313_o;
  assign n316_o = {n314_o, n305_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:990:4  */
  always @*
    case (n316_o)
      2'b10: n317_o = n309_o;
      2'b01: n317_o = n300_o;
      default: n317_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:996:12  */
  assign n318_o = q14[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:997:18  */
  assign n319_o = betaw14 - absq14d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:997:28  */
  assign n321_o = n318_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:998:18  */
  assign n322_o = betaw14 + absq14d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:996:4  */
  always @*
    case (n321_o)
      1'b1: n323_o = n319_o;
      default: n323_o = n322_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1000:18  */
  assign n324_o = w13[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1000:32  */
  assign n326_o = {n324_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1001:20  */
  assign n327_o = betaw13[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1001:38  */
  assign n328_o = d[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1001:35  */
  assign n329_o = {n327_o, n328_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1004:23  */
  assign selfunctiontable13_n330 = selfunctiontable13_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1002:4  */
  selfunction_f300_uid4 selfunctiontable13 (
    .x(sel13),
    .y(selfunctiontable13_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1009:16  */
  assign n334_o = {3'b000, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1009:66  */
  assign n336_o = q13 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1009:77  */
  assign n338_o = q13 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1009:77  */
  assign n339_o = n336_o | n338_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1010:15  */
  assign n341_o = {2'b00, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1010:22  */
  assign n343_o = {n341_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1010:52  */
  assign n345_o = q13 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1010:63  */
  assign n347_o = q13 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1010:63  */
  assign n348_o = n345_o | n347_o;
  assign n350_o = {n348_o, n339_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1007:4  */
  always @*
    case (n350_o)
      2'b10: n351_o = n343_o;
      2'b01: n351_o = n334_o;
      default: n351_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1013:12  */
  assign n352_o = q13[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1014:21  */
  assign n353_o = betaw13_d1 - absq13d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1014:31  */
  assign n355_o = n352_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1015:21  */
  assign n356_o = betaw13_d1 + absq13d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1013:4  */
  always @*
    case (n355_o)
      1'b1: n357_o = n353_o;
      default: n357_o = n356_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1017:18  */
  assign n358_o = w12[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1017:32  */
  assign n360_o = {n358_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1018:20  */
  assign n361_o = betaw12[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1018:41  */
  assign n362_o = d_d1[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1018:35  */
  assign n363_o = {n361_o, n362_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1021:23  */
  assign selfunctiontable12_n364 = selfunctiontable12_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1019:4  */
  selfunction_f300_uid4 selfunctiontable12 (
    .x(sel12),
    .y(selfunctiontable12_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1026:16  */
  assign n368_o = {3'b000, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1026:66  */
  assign n370_o = q12 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1026:77  */
  assign n372_o = q12 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1026:77  */
  assign n373_o = n370_o | n372_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1027:15  */
  assign n375_o = {2'b00, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1027:22  */
  assign n377_o = {n375_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1027:52  */
  assign n379_o = q12 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1027:63  */
  assign n381_o = q12 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1027:63  */
  assign n382_o = n379_o | n381_o;
  assign n384_o = {n382_o, n373_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1024:4  */
  always @*
    case (n384_o)
      2'b10: n385_o = n377_o;
      2'b01: n385_o = n368_o;
      default: n385_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1030:12  */
  assign n386_o = q12[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1031:21  */
  assign n387_o = betaw12_d1 - absq12d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1031:31  */
  assign n389_o = n386_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1032:21  */
  assign n390_o = betaw12_d1 + absq12d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1030:4  */
  always @*
    case (n389_o)
      1'b1: n391_o = n387_o;
      default: n391_o = n390_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1034:18  */
  assign n392_o = w11[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1034:32  */
  assign n394_o = {n392_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1035:20  */
  assign n395_o = betaw11[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1035:41  */
  assign n396_o = d_d2[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1035:35  */
  assign n397_o = {n395_o, n396_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1038:23  */
  assign selfunctiontable11_n398 = selfunctiontable11_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1036:4  */
  selfunction_f300_uid4 selfunctiontable11 (
    .x(sel11),
    .y(selfunctiontable11_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1043:16  */
  assign n402_o = {3'b000, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1043:66  */
  assign n404_o = q11 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1043:77  */
  assign n406_o = q11 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1043:77  */
  assign n407_o = n404_o | n406_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1044:15  */
  assign n409_o = {2'b00, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1044:22  */
  assign n411_o = {n409_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1044:52  */
  assign n413_o = q11 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1044:63  */
  assign n415_o = q11 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1044:63  */
  assign n416_o = n413_o | n415_o;
  assign n418_o = {n416_o, n407_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1041:4  */
  always @*
    case (n418_o)
      2'b10: n419_o = n411_o;
      2'b01: n419_o = n402_o;
      default: n419_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1047:12  */
  assign n420_o = q11[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1048:21  */
  assign n421_o = betaw11_d1 - absq11d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1048:31  */
  assign n423_o = n420_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1049:21  */
  assign n424_o = betaw11_d1 + absq11d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1047:4  */
  always @*
    case (n423_o)
      1'b1: n425_o = n421_o;
      default: n425_o = n424_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1051:18  */
  assign n426_o = w10[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1051:32  */
  assign n428_o = {n426_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1052:20  */
  assign n429_o = betaw10[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1052:41  */
  assign n430_o = d_d3[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1052:35  */
  assign n431_o = {n429_o, n430_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1055:23  */
  assign selfunctiontable10_n432 = selfunctiontable10_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1053:4  */
  selfunction_f300_uid4 selfunctiontable10 (
    .x(sel10),
    .y(selfunctiontable10_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1060:16  */
  assign n436_o = {3'b000, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1060:66  */
  assign n438_o = q10 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1060:77  */
  assign n440_o = q10 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1060:77  */
  assign n441_o = n438_o | n440_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1061:15  */
  assign n443_o = {2'b00, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1061:22  */
  assign n445_o = {n443_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1061:52  */
  assign n447_o = q10 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1061:63  */
  assign n449_o = q10 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1061:63  */
  assign n450_o = n447_o | n449_o;
  assign n452_o = {n450_o, n441_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1058:4  */
  always @*
    case (n452_o)
      2'b10: n453_o = n445_o;
      2'b01: n453_o = n436_o;
      default: n453_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1064:15  */
  assign n454_o = q10_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1065:20  */
  assign n455_o = betaw10_d1 - absq10d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1065:33  */
  assign n457_o = n454_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1066:21  */
  assign n458_o = betaw10_d1 + absq10d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1064:4  */
  always @*
    case (n457_o)
      1'b1: n459_o = n455_o;
      default: n459_o = n458_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1068:16  */
  assign n460_o = w9[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1068:30  */
  assign n462_o = {n460_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1069:18  */
  assign n463_o = betaw9[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1069:39  */
  assign n464_o = d_d4[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1069:33  */
  assign n465_o = {n463_o, n464_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1072:23  */
  assign selfunctiontable9_n466 = selfunctiontable9_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1070:4  */
  selfunction_f300_uid4 selfunctiontable9 (
    .x(sel9),
    .y(selfunctiontable9_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1077:16  */
  assign n470_o = {3'b000, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1077:66  */
  assign n472_o = q9 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1077:77  */
  assign n474_o = q9 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1077:77  */
  assign n475_o = n472_o | n474_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1078:15  */
  assign n477_o = {2'b00, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1078:22  */
  assign n479_o = {n477_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1078:52  */
  assign n481_o = q9 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1078:63  */
  assign n483_o = q9 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1078:63  */
  assign n484_o = n481_o | n483_o;
  assign n486_o = {n484_o, n475_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1075:4  */
  always @*
    case (n486_o)
      2'b10: n487_o = n479_o;
      2'b01: n487_o = n470_o;
      default: n487_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1081:14  */
  assign n488_o = q9_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1082:19  */
  assign n489_o = betaw9_d1 - absq9d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1082:31  */
  assign n491_o = n488_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1083:20  */
  assign n492_o = betaw9_d1 + absq9d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1081:4  */
  always @*
    case (n491_o)
      1'b1: n493_o = n489_o;
      default: n493_o = n492_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1085:16  */
  assign n494_o = w8[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1085:30  */
  assign n496_o = {n494_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1086:18  */
  assign n497_o = betaw8[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1086:39  */
  assign n498_o = d_d5[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1086:33  */
  assign n499_o = {n497_o, n498_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1089:23  */
  assign selfunctiontable8_n500 = selfunctiontable8_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1087:4  */
  selfunction_f300_uid4 selfunctiontable8 (
    .x(sel8),
    .y(selfunctiontable8_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1094:16  */
  assign n504_o = {3'b000, d_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1094:66  */
  assign n506_o = q8 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1094:77  */
  assign n508_o = q8 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1094:77  */
  assign n509_o = n506_o | n508_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1095:15  */
  assign n511_o = {2'b00, d_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1095:22  */
  assign n513_o = {n511_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1095:52  */
  assign n515_o = q8 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1095:63  */
  assign n517_o = q8 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1095:63  */
  assign n518_o = n515_o | n517_o;
  assign n520_o = {n518_o, n509_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1092:4  */
  always @*
    case (n520_o)
      2'b10: n521_o = n513_o;
      2'b01: n521_o = n504_o;
      default: n521_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1098:14  */
  assign n522_o = q8_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1099:19  */
  assign n523_o = betaw8_d1 - absq8d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1099:31  */
  assign n525_o = n522_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1100:20  */
  assign n526_o = betaw8_d1 + absq8d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1098:4  */
  always @*
    case (n525_o)
      1'b1: n527_o = n523_o;
      default: n527_o = n526_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1102:16  */
  assign n528_o = w7[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1102:30  */
  assign n530_o = {n528_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1103:18  */
  assign n531_o = betaw7[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1103:39  */
  assign n532_o = d_d6[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1103:33  */
  assign n533_o = {n531_o, n532_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1106:23  */
  assign selfunctiontable7_n534 = selfunctiontable7_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1104:4  */
  selfunction_f300_uid4 selfunctiontable7 (
    .x(sel7),
    .y(selfunctiontable7_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1111:16  */
  assign n538_o = {3'b000, d_d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1111:66  */
  assign n540_o = q7 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1111:77  */
  assign n542_o = q7 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1111:77  */
  assign n543_o = n540_o | n542_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1112:15  */
  assign n545_o = {2'b00, d_d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1112:22  */
  assign n547_o = {n545_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1112:52  */
  assign n549_o = q7 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1112:63  */
  assign n551_o = q7 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1112:63  */
  assign n552_o = n549_o | n551_o;
  assign n554_o = {n552_o, n543_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1109:4  */
  always @*
    case (n554_o)
      2'b10: n555_o = n547_o;
      2'b01: n555_o = n538_o;
      default: n555_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1115:11  */
  assign n556_o = q7[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1116:16  */
  assign n557_o = betaw7 - absq7d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1116:25  */
  assign n559_o = n556_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1117:17  */
  assign n560_o = betaw7 + absq7d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1115:4  */
  always @*
    case (n559_o)
      1'b1: n561_o = n557_o;
      default: n561_o = n560_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1119:16  */
  assign n562_o = w6[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1119:30  */
  assign n564_o = {n562_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1120:18  */
  assign n565_o = betaw6[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1120:39  */
  assign n566_o = d_d6[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1120:33  */
  assign n567_o = {n565_o, n566_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1123:23  */
  assign selfunctiontable6_n568 = selfunctiontable6_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1121:4  */
  selfunction_f300_uid4 selfunctiontable6 (
    .x(sel6),
    .y(selfunctiontable6_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1128:16  */
  assign n572_o = {3'b000, d_d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1128:66  */
  assign n574_o = q6 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1128:77  */
  assign n576_o = q6 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1128:77  */
  assign n577_o = n574_o | n576_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1129:15  */
  assign n579_o = {2'b00, d_d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1129:22  */
  assign n581_o = {n579_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1129:52  */
  assign n583_o = q6 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1129:63  */
  assign n585_o = q6 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1129:63  */
  assign n586_o = n583_o | n585_o;
  assign n588_o = {n586_o, n577_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1126:4  */
  always @*
    case (n588_o)
      2'b10: n589_o = n581_o;
      2'b01: n589_o = n572_o;
      default: n589_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1132:11  */
  assign n590_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1133:19  */
  assign n591_o = betaw6_d1 - absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1133:28  */
  assign n593_o = n590_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1134:20  */
  assign n594_o = betaw6_d1 + absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1132:4  */
  always @*
    case (n593_o)
      1'b1: n595_o = n591_o;
      default: n595_o = n594_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1136:16  */
  assign n596_o = w5[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1136:30  */
  assign n598_o = {n596_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1137:18  */
  assign n599_o = betaw5[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1137:39  */
  assign n600_o = d_d7[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1137:33  */
  assign n601_o = {n599_o, n600_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1140:23  */
  assign selfunctiontable5_n602 = selfunctiontable5_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1138:4  */
  selfunction_f300_uid4 selfunctiontable5 (
    .x(sel5),
    .y(selfunctiontable5_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1145:16  */
  assign n606_o = {3'b000, d_d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1145:66  */
  assign n608_o = q5 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1145:77  */
  assign n610_o = q5 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1145:77  */
  assign n611_o = n608_o | n610_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1146:15  */
  assign n613_o = {2'b00, d_d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1146:22  */
  assign n615_o = {n613_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1146:52  */
  assign n617_o = q5 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1146:63  */
  assign n619_o = q5 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1146:63  */
  assign n620_o = n617_o | n619_o;
  assign n622_o = {n620_o, n611_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1143:4  */
  always @*
    case (n622_o)
      2'b10: n623_o = n615_o;
      2'b01: n623_o = n606_o;
      default: n623_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1149:11  */
  assign n624_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1150:19  */
  assign n625_o = betaw5_d1 - absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1150:28  */
  assign n627_o = n624_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1151:20  */
  assign n628_o = betaw5_d1 + absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1149:4  */
  always @*
    case (n627_o)
      1'b1: n629_o = n625_o;
      default: n629_o = n628_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1153:16  */
  assign n630_o = w4[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1153:30  */
  assign n632_o = {n630_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1154:18  */
  assign n633_o = betaw4[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1154:39  */
  assign n634_o = d_d8[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1154:33  */
  assign n635_o = {n633_o, n634_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1157:23  */
  assign selfunctiontable4_n636 = selfunctiontable4_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1155:4  */
  selfunction_f300_uid4 selfunctiontable4 (
    .x(sel4),
    .y(selfunctiontable4_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1162:16  */
  assign n640_o = {3'b000, d_d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1162:66  */
  assign n642_o = q4 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1162:77  */
  assign n644_o = q4 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1162:77  */
  assign n645_o = n642_o | n644_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1163:15  */
  assign n647_o = {2'b00, d_d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1163:22  */
  assign n649_o = {n647_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1163:52  */
  assign n651_o = q4 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1163:63  */
  assign n653_o = q4 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1163:63  */
  assign n654_o = n651_o | n653_o;
  assign n656_o = {n654_o, n645_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1160:4  */
  always @*
    case (n656_o)
      2'b10: n657_o = n649_o;
      2'b01: n657_o = n640_o;
      default: n657_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1166:11  */
  assign n658_o = q4[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1167:19  */
  assign n659_o = betaw4_d1 - absq4d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1167:28  */
  assign n661_o = n658_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1168:20  */
  assign n662_o = betaw4_d1 + absq4d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1166:4  */
  always @*
    case (n661_o)
      1'b1: n663_o = n659_o;
      default: n663_o = n662_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1170:16  */
  assign n664_o = w3[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1170:30  */
  assign n666_o = {n664_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1171:18  */
  assign n667_o = betaw3[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1171:39  */
  assign n668_o = d_d9[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1171:33  */
  assign n669_o = {n667_o, n668_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1174:23  */
  assign selfunctiontable3_n670 = selfunctiontable3_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1172:4  */
  selfunction_f300_uid4 selfunctiontable3 (
    .x(sel3),
    .y(selfunctiontable3_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1179:16  */
  assign n674_o = {3'b000, d_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1179:66  */
  assign n676_o = q3 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1179:77  */
  assign n678_o = q3 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1179:77  */
  assign n679_o = n676_o | n678_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1180:15  */
  assign n681_o = {2'b00, d_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1180:23  */
  assign n683_o = {n681_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1180:52  */
  assign n685_o = q3 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1180:63  */
  assign n687_o = q3 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1180:63  */
  assign n688_o = n685_o | n687_o;
  assign n690_o = {n688_o, n679_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1177:4  */
  always @*
    case (n690_o)
      2'b10: n691_o = n683_o;
      2'b01: n691_o = n674_o;
      default: n691_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1183:11  */
  assign n692_o = q3[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1184:19  */
  assign n693_o = betaw3_d1 - absq3d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1184:28  */
  assign n695_o = n692_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1185:20  */
  assign n696_o = betaw3_d1 + absq3d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1183:4  */
  always @*
    case (n695_o)
      1'b1: n697_o = n693_o;
      default: n697_o = n696_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1187:16  */
  assign n698_o = w2[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1187:30  */
  assign n700_o = {n698_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1188:18  */
  assign n701_o = betaw2[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1188:40  */
  assign n702_o = d_d10[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1188:33  */
  assign n703_o = {n701_o, n702_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1191:23  */
  assign selfunctiontable2_n704 = selfunctiontable2_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1189:4  */
  selfunction_f300_uid4 selfunctiontable2 (
    .x(sel2),
    .y(selfunctiontable2_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1196:16  */
  assign n708_o = {3'b000, d_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1196:66  */
  assign n710_o = q2 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1196:77  */
  assign n712_o = q2 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1196:77  */
  assign n713_o = n710_o | n712_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1197:15  */
  assign n715_o = {2'b00, d_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1197:23  */
  assign n717_o = {n715_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1197:52  */
  assign n719_o = q2 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1197:63  */
  assign n721_o = q2 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1197:63  */
  assign n722_o = n719_o | n721_o;
  assign n724_o = {n722_o, n713_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1194:4  */
  always @*
    case (n724_o)
      2'b10: n725_o = n717_o;
      2'b01: n725_o = n708_o;
      default: n725_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1200:14  */
  assign n726_o = q2_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1201:19  */
  assign n727_o = betaw2_d1 - absq2d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1201:31  */
  assign n729_o = n726_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1202:20  */
  assign n730_o = betaw2_d1 + absq2d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1200:4  */
  always @*
    case (n729_o)
      1'b1: n731_o = n727_o;
      default: n731_o = n730_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1204:16  */
  assign n732_o = w1[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1204:30  */
  assign n734_o = {n732_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1205:18  */
  assign n735_o = betaw1[26:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1205:40  */
  assign n736_o = d_d11[22:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1205:33  */
  assign n737_o = {n735_o, n736_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1208:23  */
  assign selfunctiontable1_n738 = selfunctiontable1_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1206:4  */
  selfunction_f300_uid4 selfunctiontable1 (
    .x(sel1),
    .y(selfunctiontable1_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1213:16  */
  assign n742_o = {3'b000, d_d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1213:66  */
  assign n744_o = q1 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1213:77  */
  assign n746_o = q1 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1213:77  */
  assign n747_o = n744_o | n746_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1214:15  */
  assign n749_o = {2'b00, d_d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1214:23  */
  assign n751_o = {n749_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1214:52  */
  assign n753_o = q1 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1214:63  */
  assign n755_o = q1 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1214:63  */
  assign n756_o = n753_o | n755_o;
  assign n758_o = {n756_o, n747_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1211:4  */
  always @*
    case (n758_o)
      2'b10: n759_o = n751_o;
      2'b01: n759_o = n742_o;
      default: n759_o = 27'b000000000000000000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1217:14  */
  assign n760_o = q1_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1218:19  */
  assign n761_o = betaw1_d1 - absq1d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1218:31  */
  assign n763_o = n760_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1219:20  */
  assign n764_o = betaw1_d1 + absq1d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1217:4  */
  always @*
    case (n763_o)
      1'b1: n765_o = n761_o;
      default: n765_o = n764_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1221:16  */
  assign n766_o = w0[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1222:17  */
  assign n767_o = wfinal[24];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1223:20  */
  assign n768_o = q14[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1224:20  */
  assign n769_o = q14[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1224:24  */
  assign n771_o = {n769_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1225:20  */
  assign n772_o = q13[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1226:20  */
  assign n773_o = q13[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1226:24  */
  assign n775_o = {n773_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1227:20  */
  assign n776_o = q12[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1228:20  */
  assign n777_o = q12[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1228:24  */
  assign n779_o = {n777_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1229:20  */
  assign n780_o = q11[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1230:20  */
  assign n781_o = q11[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1230:24  */
  assign n783_o = {n781_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1231:20  */
  assign n784_o = q10[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1232:20  */
  assign n785_o = q10[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1232:24  */
  assign n787_o = {n785_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1233:18  */
  assign n788_o = q9[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1234:18  */
  assign n789_o = q9[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1234:22  */
  assign n791_o = {n789_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1235:18  */
  assign n792_o = q8[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1236:18  */
  assign n793_o = q8[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1236:22  */
  assign n795_o = {n793_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1237:18  */
  assign n796_o = q7[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1238:18  */
  assign n797_o = q7[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1238:22  */
  assign n799_o = {n797_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1239:18  */
  assign n800_o = q6[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1240:18  */
  assign n801_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1240:22  */
  assign n803_o = {n801_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1241:18  */
  assign n804_o = q5[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1242:18  */
  assign n805_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1242:22  */
  assign n807_o = {n805_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1243:18  */
  assign n808_o = q4[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1244:18  */
  assign n809_o = q4[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1244:22  */
  assign n811_o = {n809_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1245:18  */
  assign n812_o = q3[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1246:18  */
  assign n813_o = q3[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1246:22  */
  assign n815_o = {n813_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1247:18  */
  assign n816_o = q2[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1248:18  */
  assign n817_o = q2[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1248:22  */
  assign n819_o = {n817_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1249:18  */
  assign n820_o = q1[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1250:18  */
  assign n821_o = q1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1250:22  */
  assign n823_o = {n821_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:19  */
  assign n824_o = {qp14_d11, qp13_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:30  */
  assign n825_o = {n824_o, qp12_d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:40  */
  assign n826_o = {n825_o, qp11_d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:50  */
  assign n827_o = {n826_o, qp10_d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:60  */
  assign n828_o = {n827_o, qp9_d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:69  */
  assign n829_o = {n828_o, qp8_d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:78  */
  assign n830_o = {n829_o, qp7_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:87  */
  assign n831_o = {n830_o, qp6_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:96  */
  assign n832_o = {n831_o, qp5_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:105  */
  assign n833_o = {n832_o, qp4_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:114  */
  assign n834_o = {n833_o, qp3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:123  */
  assign n835_o = {n834_o, qp2_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1251:132  */
  assign n836_o = {n835_o, qp1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:18  */
  assign n837_o = qm14_d12[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:22  */
  assign n838_o = {n837_o, qm13_d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:33  */
  assign n839_o = {n838_o, qm12_d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:44  */
  assign n840_o = {n839_o, qm11_d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:54  */
  assign n841_o = {n840_o, qm10_d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:64  */
  assign n842_o = {n841_o, qm9_d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:73  */
  assign n843_o = {n842_o, qm8_d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:82  */
  assign n844_o = {n843_o, qm7_d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:91  */
  assign n845_o = {n844_o, qm6_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:100  */
  assign n846_o = {n845_o, qm5_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:109  */
  assign n847_o = {n846_o, qm4_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:118  */
  assign n848_o = {n847_o, qm3_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:127  */
  assign n849_o = {n848_o, qm2_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:136  */
  assign n850_o = {n849_o, qm1_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1252:145  */
  assign n851_o = {n850_o, qm0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1253:22  */
  assign n852_o = qp_d1 - qm;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1257:18  */
  assign n853_o = quotient[26:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1259:19  */
  assign n854_o = mr[24:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1259:41  */
  assign n855_o = mr[25];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1259:34  */
  assign n856_o = n855_o ? n854_o : n857_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1260:19  */
  assign n857_o = mr[23:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1261:19  */
  assign n858_o = frnorm[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1262:58  */
  assign n859_o = mr[25];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1262:54  */
  assign n861_o = {9'b000111111, n859_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1262:23  */
  assign n862_o = expr0_d12 + n861_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1264:29  */
  assign n863_o = frnorm[23:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1264:21  */
  assign n864_o = {expr1, n863_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1265:48  */
  assign n866_o = {32'b00000000000000000000000000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1265:24  */
  assign n867_o = expfrac + n866_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1266:36  */
  assign n869_o = expfracr[32];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1266:23  */
  assign n870_o = n869_o ? 2'b00 : n875_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1267:37  */
  assign n872_o = expfracr[32:31];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1267:52  */
  assign n874_o = n872_o == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1267:12  */
  assign n875_o = n874_o ? 2'b10 : 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1271:17  */
  assign n878_o = exnr0_d12 == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1269:4  */
  always @*
    case (n878_o)
      1'b1: n879_o = exnr;
      default: n879_o = exnr0_d12;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1273:19  */
  assign n880_o = {exnrfinal, sr_d12};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1273:38  */
  assign n881_o = expfracr[30:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:1273:28  */
  assign n882_o = {n880_o, n881_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n883_q <= expr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n884_q <= expr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n885_q <= expr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n886_q <= expr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n887_q <= expr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n888_q <= expr0_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n889_q <= expr0_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n890_q <= expr0_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n891_q <= expr0_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n892_q <= expr0_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n893_q <= expr0_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n894_q <= expr0_d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n895_q <= sr;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n896_q <= sr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n897_q <= sr_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n898_q <= sr_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n899_q <= sr_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n900_q <= sr_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n901_q <= sr_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n902_q <= sr_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n903_q <= sr_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n904_q <= sr_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n905_q <= sr_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n906_q <= sr_d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n907_q <= exnr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n908_q <= exnr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n909_q <= exnr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n910_q <= exnr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n911_q <= exnr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n912_q <= exnr0_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n913_q <= exnr0_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n914_q <= exnr0_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n915_q <= exnr0_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n916_q <= exnr0_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n917_q <= exnr0_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n918_q <= exnr0_d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n919_q <= d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n920_q <= d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n921_q <= d_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n922_q <= d_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n923_q <= d_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n924_q <= d_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n925_q <= d_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n926_q <= d_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n927_q <= d_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n928_q <= d_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n929_q <= d_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n930_q <= betaw13;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n931_q <= q13_copy6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n932_q <= betaw12;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n933_q <= q12_copy7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n934_q <= betaw11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n935_q <= q11_copy8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n936_q <= betaw10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n937_q <= q10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n938_q <= absq10d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n939_q <= betaw9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n940_q <= q9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n941_q <= absq9d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n942_q <= betaw8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n943_q <= q8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n944_q <= absq8d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n945_q <= betaw6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n946_q <= q6_copy13;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n947_q <= betaw5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n948_q <= q5_copy14;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n949_q <= betaw4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n950_q <= q4_copy15;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n951_q <= betaw3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n952_q <= q3_copy16;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n953_q <= betaw2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n954_q <= q2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n955_q <= absq2d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n956_q <= betaw1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n957_q <= q1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n958_q <= absq1d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n959_q <= qp14;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n960_q <= qp14_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n961_q <= qp14_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n962_q <= qp14_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n963_q <= qp14_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n964_q <= qp14_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n965_q <= qp14_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n966_q <= qp14_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n967_q <= qp14_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n968_q <= qp14_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n969_q <= qp14_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n970_q <= qm14;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n971_q <= qm14_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n972_q <= qm14_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n973_q <= qm14_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n974_q <= qm14_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n975_q <= qm14_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n976_q <= qm14_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n977_q <= qm14_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n978_q <= qm14_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n979_q <= qm14_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n980_q <= qm14_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n981_q <= qm14_d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n982_q <= qp13;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n983_q <= qp13_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n984_q <= qp13_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n985_q <= qp13_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n986_q <= qp13_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n987_q <= qp13_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n988_q <= qp13_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n989_q <= qp13_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n990_q <= qp13_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n991_q <= qp13_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n992_q <= qm13;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n993_q <= qm13_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n994_q <= qm13_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n995_q <= qm13_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n996_q <= qm13_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n997_q <= qm13_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n998_q <= qm13_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n999_q <= qm13_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1000_q <= qm13_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1001_q <= qm13_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1002_q <= qm13_d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1003_q <= qp12;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1004_q <= qp12_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1005_q <= qp12_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1006_q <= qp12_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1007_q <= qp12_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1008_q <= qp12_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1009_q <= qp12_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1010_q <= qp12_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1011_q <= qp12_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1012_q <= qm12;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1013_q <= qm12_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1014_q <= qm12_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1015_q <= qm12_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1016_q <= qm12_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1017_q <= qm12_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1018_q <= qm12_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1019_q <= qm12_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1020_q <= qm12_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1021_q <= qm12_d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1022_q <= qp11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1023_q <= qp11_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1024_q <= qp11_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1025_q <= qp11_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1026_q <= qp11_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1027_q <= qp11_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1028_q <= qp11_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1029_q <= qp11_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1030_q <= qm11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1031_q <= qm11_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1032_q <= qm11_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1033_q <= qm11_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1034_q <= qm11_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1035_q <= qm11_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1036_q <= qm11_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1037_q <= qm11_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1038_q <= qm11_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1039_q <= qp10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1040_q <= qp10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1041_q <= qp10_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1042_q <= qp10_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1043_q <= qp10_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1044_q <= qp10_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1045_q <= qp10_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1046_q <= qp10_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1047_q <= qm10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1048_q <= qm10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1049_q <= qm10_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1050_q <= qm10_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1051_q <= qm10_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1052_q <= qm10_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1053_q <= qm10_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1054_q <= qm10_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1055_q <= qm10_d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1056_q <= qp9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1057_q <= qp9_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1058_q <= qp9_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1059_q <= qp9_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1060_q <= qp9_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1061_q <= qp9_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1062_q <= qp9_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1063_q <= qm9;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1064_q <= qm9_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1065_q <= qm9_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1066_q <= qm9_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1067_q <= qm9_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1068_q <= qm9_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1069_q <= qm9_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1070_q <= qm9_d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1071_q <= qp8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1072_q <= qp8_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1073_q <= qp8_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1074_q <= qp8_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1075_q <= qp8_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1076_q <= qp8_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1077_q <= qm8;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1078_q <= qm8_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1079_q <= qm8_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1080_q <= qm8_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1081_q <= qm8_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1082_q <= qm8_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1083_q <= qm8_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1084_q <= qp7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1085_q <= qp7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1086_q <= qp7_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1087_q <= qp7_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1088_q <= qp7_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1089_q <= qm7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1090_q <= qm7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1091_q <= qm7_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1092_q <= qm7_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1093_q <= qm7_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1094_q <= qm7_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1095_q <= qp6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1096_q <= qp6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1097_q <= qp6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1098_q <= qp6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1099_q <= qm6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1100_q <= qm6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1101_q <= qm6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1102_q <= qm6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1103_q <= qm6_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1104_q <= qp5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1105_q <= qp5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1106_q <= qp5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1107_q <= qm5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1108_q <= qm5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1109_q <= qm5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1110_q <= qm5_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1111_q <= qp4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1112_q <= qp4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1113_q <= qm4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1114_q <= qm4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1115_q <= qm4_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1116_q <= qp3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1117_q <= qm3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1118_q <= qm3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1119_q <= qp2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1120_q <= qm2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1121_q <= qm2_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1122_q <= qm1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_8_23.vhdl:724:10  */
  always @(posedge clk)
    n1123_q <= qp;
endmodule

