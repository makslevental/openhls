module selfunction_f300_uid4
  (input wire [8:0] x,
   output wire [2:0] y);
  wire [2:0] y0;
  wire [2:0] y1;
  wire n433_o;
  wire n436_o;
  wire n439_o;
  wire n442_o;
  wire n445_o;
  wire n448_o;
  wire n451_o;
  wire n454_o;
  wire n457_o;
  wire n460_o;
  wire n463_o;
  wire n466_o;
  wire n469_o;
  wire n472_o;
  wire n475_o;
  wire n478_o;
  wire n481_o;
  wire n484_o;
  wire n487_o;
  wire n490_o;
  wire n493_o;
  wire n496_o;
  wire n499_o;
  wire n502_o;
  wire n505_o;
  wire n508_o;
  wire n511_o;
  wire n514_o;
  wire n517_o;
  wire n520_o;
  wire n523_o;
  wire n526_o;
  wire n529_o;
  wire n532_o;
  wire n535_o;
  wire n538_o;
  wire n541_o;
  wire n544_o;
  wire n547_o;
  wire n550_o;
  wire n553_o;
  wire n556_o;
  wire n559_o;
  wire n562_o;
  wire n565_o;
  wire n568_o;
  wire n571_o;
  wire n574_o;
  wire n577_o;
  wire n580_o;
  wire n583_o;
  wire n586_o;
  wire n589_o;
  wire n592_o;
  wire n595_o;
  wire n598_o;
  wire n601_o;
  wire n604_o;
  wire n607_o;
  wire n610_o;
  wire n613_o;
  wire n616_o;
  wire n619_o;
  wire n622_o;
  wire n625_o;
  wire n628_o;
  wire n631_o;
  wire n634_o;
  wire n637_o;
  wire n640_o;
  wire n643_o;
  wire n646_o;
  wire n649_o;
  wire n652_o;
  wire n655_o;
  wire n658_o;
  wire n661_o;
  wire n664_o;
  wire n667_o;
  wire n670_o;
  wire n673_o;
  wire n676_o;
  wire n679_o;
  wire n682_o;
  wire n685_o;
  wire n688_o;
  wire n691_o;
  wire n694_o;
  wire n697_o;
  wire n700_o;
  wire n703_o;
  wire n706_o;
  wire n709_o;
  wire n712_o;
  wire n715_o;
  wire n718_o;
  wire n721_o;
  wire n724_o;
  wire n727_o;
  wire n730_o;
  wire n733_o;
  wire n736_o;
  wire n739_o;
  wire n742_o;
  wire n745_o;
  wire n748_o;
  wire n751_o;
  wire n754_o;
  wire n757_o;
  wire n760_o;
  wire n763_o;
  wire n766_o;
  wire n769_o;
  wire n772_o;
  wire n775_o;
  wire n778_o;
  wire n781_o;
  wire n784_o;
  wire n787_o;
  wire n790_o;
  wire n793_o;
  wire n796_o;
  wire n799_o;
  wire n802_o;
  wire n805_o;
  wire n808_o;
  wire n811_o;
  wire n814_o;
  wire n817_o;
  wire n820_o;
  wire n823_o;
  wire n826_o;
  wire n829_o;
  wire n832_o;
  wire n835_o;
  wire n838_o;
  wire n841_o;
  wire n844_o;
  wire n847_o;
  wire n850_o;
  wire n853_o;
  wire n856_o;
  wire n859_o;
  wire n862_o;
  wire n865_o;
  wire n868_o;
  wire n871_o;
  wire n874_o;
  wire n877_o;
  wire n880_o;
  wire n883_o;
  wire n886_o;
  wire n889_o;
  wire n892_o;
  wire n895_o;
  wire n898_o;
  wire n901_o;
  wire n904_o;
  wire n907_o;
  wire n910_o;
  wire n913_o;
  wire n916_o;
  wire n919_o;
  wire n922_o;
  wire n925_o;
  wire n928_o;
  wire n931_o;
  wire n934_o;
  wire n937_o;
  wire n940_o;
  wire n943_o;
  wire n946_o;
  wire n949_o;
  wire n952_o;
  wire n955_o;
  wire n958_o;
  wire n961_o;
  wire n964_o;
  wire n967_o;
  wire n970_o;
  wire n973_o;
  wire n976_o;
  wire n979_o;
  wire n982_o;
  wire n985_o;
  wire n988_o;
  wire n991_o;
  wire n994_o;
  wire n997_o;
  wire n1000_o;
  wire n1003_o;
  wire n1006_o;
  wire n1009_o;
  wire n1012_o;
  wire n1015_o;
  wire n1018_o;
  wire n1021_o;
  wire n1024_o;
  wire n1027_o;
  wire n1030_o;
  wire n1033_o;
  wire n1036_o;
  wire n1039_o;
  wire n1042_o;
  wire n1045_o;
  wire n1048_o;
  wire n1051_o;
  wire n1054_o;
  wire n1057_o;
  wire n1060_o;
  wire n1063_o;
  wire n1066_o;
  wire n1069_o;
  wire n1072_o;
  wire n1075_o;
  wire n1078_o;
  wire n1081_o;
  wire n1084_o;
  wire n1087_o;
  wire n1090_o;
  wire n1093_o;
  wire n1096_o;
  wire n1099_o;
  wire n1102_o;
  wire n1105_o;
  wire n1108_o;
  wire n1111_o;
  wire n1114_o;
  wire n1117_o;
  wire n1120_o;
  wire n1123_o;
  wire n1126_o;
  wire n1129_o;
  wire n1132_o;
  wire n1135_o;
  wire n1138_o;
  wire n1141_o;
  wire n1144_o;
  wire n1147_o;
  wire n1150_o;
  wire n1153_o;
  wire n1156_o;
  wire n1159_o;
  wire n1162_o;
  wire n1165_o;
  wire n1168_o;
  wire n1171_o;
  wire n1174_o;
  wire n1177_o;
  wire n1180_o;
  wire n1183_o;
  wire n1186_o;
  wire n1189_o;
  wire n1192_o;
  wire n1195_o;
  wire n1198_o;
  wire n1201_o;
  wire n1204_o;
  wire n1207_o;
  wire n1210_o;
  wire n1213_o;
  wire n1216_o;
  wire n1219_o;
  wire n1222_o;
  wire n1225_o;
  wire n1228_o;
  wire n1231_o;
  wire n1234_o;
  wire n1237_o;
  wire n1240_o;
  wire n1243_o;
  wire n1246_o;
  wire n1249_o;
  wire n1252_o;
  wire n1255_o;
  wire n1258_o;
  wire n1261_o;
  wire n1264_o;
  wire n1267_o;
  wire n1270_o;
  wire n1273_o;
  wire n1276_o;
  wire n1279_o;
  wire n1282_o;
  wire n1285_o;
  wire n1288_o;
  wire n1291_o;
  wire n1294_o;
  wire n1297_o;
  wire n1300_o;
  wire n1303_o;
  wire n1306_o;
  wire n1309_o;
  wire n1312_o;
  wire n1315_o;
  wire n1318_o;
  wire n1321_o;
  wire n1324_o;
  wire n1327_o;
  wire n1330_o;
  wire n1333_o;
  wire n1336_o;
  wire n1339_o;
  wire n1342_o;
  wire n1345_o;
  wire n1348_o;
  wire n1351_o;
  wire n1354_o;
  wire n1357_o;
  wire n1360_o;
  wire n1363_o;
  wire n1366_o;
  wire n1369_o;
  wire n1372_o;
  wire n1375_o;
  wire n1378_o;
  wire n1381_o;
  wire n1384_o;
  wire n1387_o;
  wire n1390_o;
  wire n1393_o;
  wire n1396_o;
  wire n1399_o;
  wire n1402_o;
  wire n1405_o;
  wire n1408_o;
  wire n1411_o;
  wire n1414_o;
  wire n1417_o;
  wire n1420_o;
  wire n1423_o;
  wire n1426_o;
  wire n1429_o;
  wire n1432_o;
  wire n1435_o;
  wire n1438_o;
  wire n1441_o;
  wire n1444_o;
  wire n1447_o;
  wire n1450_o;
  wire n1453_o;
  wire n1456_o;
  wire n1459_o;
  wire n1462_o;
  wire n1465_o;
  wire n1468_o;
  wire n1471_o;
  wire n1474_o;
  wire n1477_o;
  wire n1480_o;
  wire n1483_o;
  wire n1486_o;
  wire n1489_o;
  wire n1492_o;
  wire n1495_o;
  wire n1498_o;
  wire n1501_o;
  wire n1504_o;
  wire n1507_o;
  wire n1510_o;
  wire n1513_o;
  wire n1516_o;
  wire n1519_o;
  wire n1522_o;
  wire n1525_o;
  wire n1528_o;
  wire n1531_o;
  wire n1534_o;
  wire n1537_o;
  wire n1540_o;
  wire n1543_o;
  wire n1546_o;
  wire n1549_o;
  wire n1552_o;
  wire n1555_o;
  wire n1558_o;
  wire n1561_o;
  wire n1564_o;
  wire n1567_o;
  wire n1570_o;
  wire n1573_o;
  wire n1576_o;
  wire n1579_o;
  wire n1582_o;
  wire n1585_o;
  wire n1588_o;
  wire n1591_o;
  wire n1594_o;
  wire n1597_o;
  wire n1600_o;
  wire n1603_o;
  wire n1606_o;
  wire n1609_o;
  wire n1612_o;
  wire n1615_o;
  wire n1618_o;
  wire n1621_o;
  wire n1624_o;
  wire n1627_o;
  wire n1630_o;
  wire n1633_o;
  wire n1636_o;
  wire n1639_o;
  wire n1642_o;
  wire n1645_o;
  wire n1648_o;
  wire n1651_o;
  wire n1654_o;
  wire n1657_o;
  wire n1660_o;
  wire n1663_o;
  wire n1666_o;
  wire n1669_o;
  wire n1672_o;
  wire n1675_o;
  wire n1678_o;
  wire n1681_o;
  wire n1684_o;
  wire n1687_o;
  wire n1690_o;
  wire n1693_o;
  wire n1696_o;
  wire n1699_o;
  wire n1702_o;
  wire n1705_o;
  wire n1708_o;
  wire n1711_o;
  wire n1714_o;
  wire n1717_o;
  wire n1720_o;
  wire n1723_o;
  wire n1726_o;
  wire n1729_o;
  wire n1732_o;
  wire n1735_o;
  wire n1738_o;
  wire n1741_o;
  wire n1744_o;
  wire n1747_o;
  wire n1750_o;
  wire n1753_o;
  wire n1756_o;
  wire n1759_o;
  wire n1762_o;
  wire n1765_o;
  wire n1768_o;
  wire n1771_o;
  wire n1774_o;
  wire n1777_o;
  wire n1780_o;
  wire n1783_o;
  wire n1786_o;
  wire n1789_o;
  wire n1792_o;
  wire n1795_o;
  wire n1798_o;
  wire n1801_o;
  wire n1804_o;
  wire n1807_o;
  wire n1810_o;
  wire n1813_o;
  wire n1816_o;
  wire n1819_o;
  wire n1822_o;
  wire n1825_o;
  wire n1828_o;
  wire n1831_o;
  wire n1834_o;
  wire n1837_o;
  wire n1840_o;
  wire n1843_o;
  wire n1846_o;
  wire n1849_o;
  wire n1852_o;
  wire n1855_o;
  wire n1858_o;
  wire n1861_o;
  wire n1864_o;
  wire n1867_o;
  wire n1870_o;
  wire n1873_o;
  wire n1876_o;
  wire n1879_o;
  wire n1882_o;
  wire n1885_o;
  wire n1888_o;
  wire n1891_o;
  wire n1894_o;
  wire n1897_o;
  wire n1900_o;
  wire n1903_o;
  wire n1906_o;
  wire n1909_o;
  wire n1912_o;
  wire n1915_o;
  wire n1918_o;
  wire n1921_o;
  wire n1924_o;
  wire n1927_o;
  wire n1930_o;
  wire n1933_o;
  wire n1936_o;
  wire n1939_o;
  wire n1942_o;
  wire n1945_o;
  wire n1948_o;
  wire n1951_o;
  wire n1954_o;
  wire n1957_o;
  wire n1960_o;
  wire n1963_o;
  wire n1966_o;
  wire [511:0] n1968_o;
  reg [2:0] n1969_o;
  assign y = y1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:28:8  */
  assign y0 = n1969_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:33:8  */
  assign y1 = y0; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:36:13  */
  assign n433_o = x == 9'b000000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:37:13  */
  assign n436_o = x == 9'b000000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:38:13  */
  assign n439_o = x == 9'b000000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:39:13  */
  assign n442_o = x == 9'b000000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:40:13  */
  assign n445_o = x == 9'b000000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:41:13  */
  assign n448_o = x == 9'b000000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:42:13  */
  assign n451_o = x == 9'b000000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:43:13  */
  assign n454_o = x == 9'b000000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:44:13  */
  assign n457_o = x == 9'b000001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:45:13  */
  assign n460_o = x == 9'b000001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:46:13  */
  assign n463_o = x == 9'b000001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:47:13  */
  assign n466_o = x == 9'b000001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:48:13  */
  assign n469_o = x == 9'b000001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:49:13  */
  assign n472_o = x == 9'b000001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:50:13  */
  assign n475_o = x == 9'b000001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:51:13  */
  assign n478_o = x == 9'b000001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:52:13  */
  assign n481_o = x == 9'b000010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:53:13  */
  assign n484_o = x == 9'b000010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:54:13  */
  assign n487_o = x == 9'b000010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:55:13  */
  assign n490_o = x == 9'b000010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:56:13  */
  assign n493_o = x == 9'b000010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:57:13  */
  assign n496_o = x == 9'b000010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:58:13  */
  assign n499_o = x == 9'b000010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:59:13  */
  assign n502_o = x == 9'b000010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:60:13  */
  assign n505_o = x == 9'b000011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:61:13  */
  assign n508_o = x == 9'b000011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:62:13  */
  assign n511_o = x == 9'b000011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:63:13  */
  assign n514_o = x == 9'b000011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:64:13  */
  assign n517_o = x == 9'b000011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:65:13  */
  assign n520_o = x == 9'b000011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:66:13  */
  assign n523_o = x == 9'b000011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:67:13  */
  assign n526_o = x == 9'b000011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:68:13  */
  assign n529_o = x == 9'b000100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:69:13  */
  assign n532_o = x == 9'b000100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:70:13  */
  assign n535_o = x == 9'b000100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:71:13  */
  assign n538_o = x == 9'b000100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:72:13  */
  assign n541_o = x == 9'b000100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:73:13  */
  assign n544_o = x == 9'b000100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:74:13  */
  assign n547_o = x == 9'b000100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:75:13  */
  assign n550_o = x == 9'b000100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:76:13  */
  assign n553_o = x == 9'b000101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:77:13  */
  assign n556_o = x == 9'b000101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:78:13  */
  assign n559_o = x == 9'b000101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:79:13  */
  assign n562_o = x == 9'b000101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:80:13  */
  assign n565_o = x == 9'b000101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:81:13  */
  assign n568_o = x == 9'b000101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:82:13  */
  assign n571_o = x == 9'b000101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:83:13  */
  assign n574_o = x == 9'b000101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:84:13  */
  assign n577_o = x == 9'b000110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:85:13  */
  assign n580_o = x == 9'b000110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:86:13  */
  assign n583_o = x == 9'b000110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:87:13  */
  assign n586_o = x == 9'b000110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:88:13  */
  assign n589_o = x == 9'b000110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:89:13  */
  assign n592_o = x == 9'b000110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:90:13  */
  assign n595_o = x == 9'b000110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:91:13  */
  assign n598_o = x == 9'b000110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:92:13  */
  assign n601_o = x == 9'b000111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:93:13  */
  assign n604_o = x == 9'b000111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:94:13  */
  assign n607_o = x == 9'b000111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:95:13  */
  assign n610_o = x == 9'b000111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:96:13  */
  assign n613_o = x == 9'b000111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:97:13  */
  assign n616_o = x == 9'b000111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:98:13  */
  assign n619_o = x == 9'b000111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:99:13  */
  assign n622_o = x == 9'b000111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:100:13  */
  assign n625_o = x == 9'b001000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:101:13  */
  assign n628_o = x == 9'b001000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:102:13  */
  assign n631_o = x == 9'b001000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:103:13  */
  assign n634_o = x == 9'b001000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:104:13  */
  assign n637_o = x == 9'b001000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:105:13  */
  assign n640_o = x == 9'b001000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:106:13  */
  assign n643_o = x == 9'b001000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:107:13  */
  assign n646_o = x == 9'b001000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:108:13  */
  assign n649_o = x == 9'b001001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:109:13  */
  assign n652_o = x == 9'b001001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:110:13  */
  assign n655_o = x == 9'b001001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:111:13  */
  assign n658_o = x == 9'b001001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:112:13  */
  assign n661_o = x == 9'b001001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:113:13  */
  assign n664_o = x == 9'b001001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:114:13  */
  assign n667_o = x == 9'b001001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:115:13  */
  assign n670_o = x == 9'b001001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:116:13  */
  assign n673_o = x == 9'b001010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:117:13  */
  assign n676_o = x == 9'b001010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:118:13  */
  assign n679_o = x == 9'b001010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:119:13  */
  assign n682_o = x == 9'b001010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:120:13  */
  assign n685_o = x == 9'b001010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:121:13  */
  assign n688_o = x == 9'b001010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:122:13  */
  assign n691_o = x == 9'b001010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:123:13  */
  assign n694_o = x == 9'b001010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:124:13  */
  assign n697_o = x == 9'b001011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:125:13  */
  assign n700_o = x == 9'b001011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:126:13  */
  assign n703_o = x == 9'b001011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:127:13  */
  assign n706_o = x == 9'b001011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:128:13  */
  assign n709_o = x == 9'b001011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:129:13  */
  assign n712_o = x == 9'b001011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:130:13  */
  assign n715_o = x == 9'b001011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:131:13  */
  assign n718_o = x == 9'b001011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:132:13  */
  assign n721_o = x == 9'b001100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:133:13  */
  assign n724_o = x == 9'b001100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:134:13  */
  assign n727_o = x == 9'b001100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:135:13  */
  assign n730_o = x == 9'b001100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:136:13  */
  assign n733_o = x == 9'b001100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:137:13  */
  assign n736_o = x == 9'b001100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:138:13  */
  assign n739_o = x == 9'b001100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:139:13  */
  assign n742_o = x == 9'b001100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:140:13  */
  assign n745_o = x == 9'b001101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:141:13  */
  assign n748_o = x == 9'b001101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:142:13  */
  assign n751_o = x == 9'b001101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:143:13  */
  assign n754_o = x == 9'b001101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:144:13  */
  assign n757_o = x == 9'b001101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:145:13  */
  assign n760_o = x == 9'b001101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:146:13  */
  assign n763_o = x == 9'b001101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:147:13  */
  assign n766_o = x == 9'b001101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:148:13  */
  assign n769_o = x == 9'b001110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:149:13  */
  assign n772_o = x == 9'b001110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:150:13  */
  assign n775_o = x == 9'b001110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:151:13  */
  assign n778_o = x == 9'b001110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:152:13  */
  assign n781_o = x == 9'b001110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:153:13  */
  assign n784_o = x == 9'b001110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:154:13  */
  assign n787_o = x == 9'b001110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:155:13  */
  assign n790_o = x == 9'b001110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:156:13  */
  assign n793_o = x == 9'b001111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:157:13  */
  assign n796_o = x == 9'b001111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:158:13  */
  assign n799_o = x == 9'b001111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:159:13  */
  assign n802_o = x == 9'b001111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:160:13  */
  assign n805_o = x == 9'b001111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:161:13  */
  assign n808_o = x == 9'b001111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:162:13  */
  assign n811_o = x == 9'b001111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:163:13  */
  assign n814_o = x == 9'b001111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:164:13  */
  assign n817_o = x == 9'b010000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:165:13  */
  assign n820_o = x == 9'b010000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:166:13  */
  assign n823_o = x == 9'b010000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:167:13  */
  assign n826_o = x == 9'b010000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:168:13  */
  assign n829_o = x == 9'b010000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:169:13  */
  assign n832_o = x == 9'b010000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:170:13  */
  assign n835_o = x == 9'b010000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:171:13  */
  assign n838_o = x == 9'b010000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:172:13  */
  assign n841_o = x == 9'b010001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:173:13  */
  assign n844_o = x == 9'b010001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:174:13  */
  assign n847_o = x == 9'b010001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:175:13  */
  assign n850_o = x == 9'b010001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:176:13  */
  assign n853_o = x == 9'b010001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:177:13  */
  assign n856_o = x == 9'b010001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:178:13  */
  assign n859_o = x == 9'b010001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:179:13  */
  assign n862_o = x == 9'b010001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:180:13  */
  assign n865_o = x == 9'b010010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:181:13  */
  assign n868_o = x == 9'b010010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:182:13  */
  assign n871_o = x == 9'b010010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:183:13  */
  assign n874_o = x == 9'b010010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:184:13  */
  assign n877_o = x == 9'b010010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:185:13  */
  assign n880_o = x == 9'b010010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:186:13  */
  assign n883_o = x == 9'b010010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:187:13  */
  assign n886_o = x == 9'b010010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:188:13  */
  assign n889_o = x == 9'b010011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:189:13  */
  assign n892_o = x == 9'b010011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:190:13  */
  assign n895_o = x == 9'b010011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:191:13  */
  assign n898_o = x == 9'b010011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:192:13  */
  assign n901_o = x == 9'b010011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:193:13  */
  assign n904_o = x == 9'b010011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:194:13  */
  assign n907_o = x == 9'b010011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:195:13  */
  assign n910_o = x == 9'b010011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:196:13  */
  assign n913_o = x == 9'b010100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:197:13  */
  assign n916_o = x == 9'b010100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:198:13  */
  assign n919_o = x == 9'b010100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:199:13  */
  assign n922_o = x == 9'b010100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:200:13  */
  assign n925_o = x == 9'b010100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:201:13  */
  assign n928_o = x == 9'b010100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:202:13  */
  assign n931_o = x == 9'b010100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:203:13  */
  assign n934_o = x == 9'b010100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:204:13  */
  assign n937_o = x == 9'b010101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:205:13  */
  assign n940_o = x == 9'b010101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:206:13  */
  assign n943_o = x == 9'b010101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:207:13  */
  assign n946_o = x == 9'b010101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:208:13  */
  assign n949_o = x == 9'b010101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:209:13  */
  assign n952_o = x == 9'b010101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:210:13  */
  assign n955_o = x == 9'b010101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:211:13  */
  assign n958_o = x == 9'b010101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:212:13  */
  assign n961_o = x == 9'b010110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:213:13  */
  assign n964_o = x == 9'b010110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:214:13  */
  assign n967_o = x == 9'b010110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:215:13  */
  assign n970_o = x == 9'b010110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:216:13  */
  assign n973_o = x == 9'b010110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:217:13  */
  assign n976_o = x == 9'b010110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:218:13  */
  assign n979_o = x == 9'b010110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:219:13  */
  assign n982_o = x == 9'b010110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:220:13  */
  assign n985_o = x == 9'b010111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:221:13  */
  assign n988_o = x == 9'b010111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:222:13  */
  assign n991_o = x == 9'b010111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:223:13  */
  assign n994_o = x == 9'b010111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:224:13  */
  assign n997_o = x == 9'b010111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:225:13  */
  assign n1000_o = x == 9'b010111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:226:13  */
  assign n1003_o = x == 9'b010111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:227:13  */
  assign n1006_o = x == 9'b010111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:228:13  */
  assign n1009_o = x == 9'b011000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:229:13  */
  assign n1012_o = x == 9'b011000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:230:13  */
  assign n1015_o = x == 9'b011000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:231:13  */
  assign n1018_o = x == 9'b011000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:232:13  */
  assign n1021_o = x == 9'b011000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:233:13  */
  assign n1024_o = x == 9'b011000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:234:13  */
  assign n1027_o = x == 9'b011000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:235:13  */
  assign n1030_o = x == 9'b011000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:236:13  */
  assign n1033_o = x == 9'b011001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:237:13  */
  assign n1036_o = x == 9'b011001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:238:13  */
  assign n1039_o = x == 9'b011001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:239:13  */
  assign n1042_o = x == 9'b011001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:240:13  */
  assign n1045_o = x == 9'b011001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:241:13  */
  assign n1048_o = x == 9'b011001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:242:13  */
  assign n1051_o = x == 9'b011001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:243:13  */
  assign n1054_o = x == 9'b011001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:244:13  */
  assign n1057_o = x == 9'b011010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:245:13  */
  assign n1060_o = x == 9'b011010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:246:13  */
  assign n1063_o = x == 9'b011010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:247:13  */
  assign n1066_o = x == 9'b011010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:248:13  */
  assign n1069_o = x == 9'b011010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:249:13  */
  assign n1072_o = x == 9'b011010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:250:13  */
  assign n1075_o = x == 9'b011010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:251:13  */
  assign n1078_o = x == 9'b011010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:252:13  */
  assign n1081_o = x == 9'b011011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:253:13  */
  assign n1084_o = x == 9'b011011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:254:13  */
  assign n1087_o = x == 9'b011011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:255:13  */
  assign n1090_o = x == 9'b011011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:256:13  */
  assign n1093_o = x == 9'b011011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:257:13  */
  assign n1096_o = x == 9'b011011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:258:13  */
  assign n1099_o = x == 9'b011011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:259:13  */
  assign n1102_o = x == 9'b011011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:260:13  */
  assign n1105_o = x == 9'b011100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:261:13  */
  assign n1108_o = x == 9'b011100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:262:13  */
  assign n1111_o = x == 9'b011100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:263:13  */
  assign n1114_o = x == 9'b011100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:264:13  */
  assign n1117_o = x == 9'b011100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:265:13  */
  assign n1120_o = x == 9'b011100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:266:13  */
  assign n1123_o = x == 9'b011100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:267:13  */
  assign n1126_o = x == 9'b011100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:268:13  */
  assign n1129_o = x == 9'b011101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:269:13  */
  assign n1132_o = x == 9'b011101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:270:13  */
  assign n1135_o = x == 9'b011101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:271:13  */
  assign n1138_o = x == 9'b011101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:272:13  */
  assign n1141_o = x == 9'b011101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:273:13  */
  assign n1144_o = x == 9'b011101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:274:13  */
  assign n1147_o = x == 9'b011101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:275:13  */
  assign n1150_o = x == 9'b011101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:276:13  */
  assign n1153_o = x == 9'b011110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:277:13  */
  assign n1156_o = x == 9'b011110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:278:13  */
  assign n1159_o = x == 9'b011110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:279:13  */
  assign n1162_o = x == 9'b011110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:280:13  */
  assign n1165_o = x == 9'b011110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:281:13  */
  assign n1168_o = x == 9'b011110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:282:13  */
  assign n1171_o = x == 9'b011110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:283:13  */
  assign n1174_o = x == 9'b011110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:284:13  */
  assign n1177_o = x == 9'b011111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:285:13  */
  assign n1180_o = x == 9'b011111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:286:13  */
  assign n1183_o = x == 9'b011111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:287:13  */
  assign n1186_o = x == 9'b011111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:288:13  */
  assign n1189_o = x == 9'b011111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:289:13  */
  assign n1192_o = x == 9'b011111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:290:13  */
  assign n1195_o = x == 9'b011111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:291:13  */
  assign n1198_o = x == 9'b011111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:292:13  */
  assign n1201_o = x == 9'b100000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:293:13  */
  assign n1204_o = x == 9'b100000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:294:13  */
  assign n1207_o = x == 9'b100000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:295:13  */
  assign n1210_o = x == 9'b100000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:296:13  */
  assign n1213_o = x == 9'b100000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:297:13  */
  assign n1216_o = x == 9'b100000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:298:13  */
  assign n1219_o = x == 9'b100000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:299:13  */
  assign n1222_o = x == 9'b100000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:300:13  */
  assign n1225_o = x == 9'b100001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:301:13  */
  assign n1228_o = x == 9'b100001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:302:13  */
  assign n1231_o = x == 9'b100001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:303:13  */
  assign n1234_o = x == 9'b100001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:304:13  */
  assign n1237_o = x == 9'b100001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:305:13  */
  assign n1240_o = x == 9'b100001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:306:13  */
  assign n1243_o = x == 9'b100001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:307:13  */
  assign n1246_o = x == 9'b100001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:308:13  */
  assign n1249_o = x == 9'b100010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:309:13  */
  assign n1252_o = x == 9'b100010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:310:13  */
  assign n1255_o = x == 9'b100010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:311:13  */
  assign n1258_o = x == 9'b100010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:312:13  */
  assign n1261_o = x == 9'b100010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:313:13  */
  assign n1264_o = x == 9'b100010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:314:13  */
  assign n1267_o = x == 9'b100010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:315:13  */
  assign n1270_o = x == 9'b100010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:316:13  */
  assign n1273_o = x == 9'b100011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:317:13  */
  assign n1276_o = x == 9'b100011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:318:13  */
  assign n1279_o = x == 9'b100011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:319:13  */
  assign n1282_o = x == 9'b100011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:320:13  */
  assign n1285_o = x == 9'b100011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:321:13  */
  assign n1288_o = x == 9'b100011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:322:13  */
  assign n1291_o = x == 9'b100011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:323:13  */
  assign n1294_o = x == 9'b100011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:324:13  */
  assign n1297_o = x == 9'b100100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:325:13  */
  assign n1300_o = x == 9'b100100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:326:13  */
  assign n1303_o = x == 9'b100100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:327:13  */
  assign n1306_o = x == 9'b100100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:328:13  */
  assign n1309_o = x == 9'b100100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:329:13  */
  assign n1312_o = x == 9'b100100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:330:13  */
  assign n1315_o = x == 9'b100100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:331:13  */
  assign n1318_o = x == 9'b100100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:332:13  */
  assign n1321_o = x == 9'b100101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:333:13  */
  assign n1324_o = x == 9'b100101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:334:13  */
  assign n1327_o = x == 9'b100101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:335:13  */
  assign n1330_o = x == 9'b100101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:336:13  */
  assign n1333_o = x == 9'b100101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:337:13  */
  assign n1336_o = x == 9'b100101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:338:13  */
  assign n1339_o = x == 9'b100101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:339:13  */
  assign n1342_o = x == 9'b100101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:340:13  */
  assign n1345_o = x == 9'b100110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:341:13  */
  assign n1348_o = x == 9'b100110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:342:13  */
  assign n1351_o = x == 9'b100110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:343:13  */
  assign n1354_o = x == 9'b100110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:344:13  */
  assign n1357_o = x == 9'b100110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:345:13  */
  assign n1360_o = x == 9'b100110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:346:13  */
  assign n1363_o = x == 9'b100110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:347:13  */
  assign n1366_o = x == 9'b100110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:348:13  */
  assign n1369_o = x == 9'b100111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:349:13  */
  assign n1372_o = x == 9'b100111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:350:13  */
  assign n1375_o = x == 9'b100111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:351:13  */
  assign n1378_o = x == 9'b100111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:352:13  */
  assign n1381_o = x == 9'b100111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:353:13  */
  assign n1384_o = x == 9'b100111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:354:13  */
  assign n1387_o = x == 9'b100111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:355:13  */
  assign n1390_o = x == 9'b100111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:356:13  */
  assign n1393_o = x == 9'b101000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:357:13  */
  assign n1396_o = x == 9'b101000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:358:13  */
  assign n1399_o = x == 9'b101000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:359:13  */
  assign n1402_o = x == 9'b101000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:360:13  */
  assign n1405_o = x == 9'b101000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:361:13  */
  assign n1408_o = x == 9'b101000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:362:13  */
  assign n1411_o = x == 9'b101000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:363:13  */
  assign n1414_o = x == 9'b101000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:364:13  */
  assign n1417_o = x == 9'b101001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:365:13  */
  assign n1420_o = x == 9'b101001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:366:13  */
  assign n1423_o = x == 9'b101001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:367:13  */
  assign n1426_o = x == 9'b101001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:368:13  */
  assign n1429_o = x == 9'b101001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:369:13  */
  assign n1432_o = x == 9'b101001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:370:13  */
  assign n1435_o = x == 9'b101001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:371:13  */
  assign n1438_o = x == 9'b101001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:372:13  */
  assign n1441_o = x == 9'b101010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:373:13  */
  assign n1444_o = x == 9'b101010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:374:13  */
  assign n1447_o = x == 9'b101010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:375:13  */
  assign n1450_o = x == 9'b101010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:376:13  */
  assign n1453_o = x == 9'b101010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:377:13  */
  assign n1456_o = x == 9'b101010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:378:13  */
  assign n1459_o = x == 9'b101010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:379:13  */
  assign n1462_o = x == 9'b101010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:380:13  */
  assign n1465_o = x == 9'b101011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:381:13  */
  assign n1468_o = x == 9'b101011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:382:13  */
  assign n1471_o = x == 9'b101011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:383:13  */
  assign n1474_o = x == 9'b101011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:384:13  */
  assign n1477_o = x == 9'b101011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:385:13  */
  assign n1480_o = x == 9'b101011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:386:13  */
  assign n1483_o = x == 9'b101011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:387:13  */
  assign n1486_o = x == 9'b101011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:388:13  */
  assign n1489_o = x == 9'b101100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:389:13  */
  assign n1492_o = x == 9'b101100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:390:13  */
  assign n1495_o = x == 9'b101100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:391:13  */
  assign n1498_o = x == 9'b101100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:392:13  */
  assign n1501_o = x == 9'b101100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:393:13  */
  assign n1504_o = x == 9'b101100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:394:13  */
  assign n1507_o = x == 9'b101100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:395:13  */
  assign n1510_o = x == 9'b101100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:396:13  */
  assign n1513_o = x == 9'b101101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:397:13  */
  assign n1516_o = x == 9'b101101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:398:13  */
  assign n1519_o = x == 9'b101101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:399:13  */
  assign n1522_o = x == 9'b101101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:400:13  */
  assign n1525_o = x == 9'b101101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:401:13  */
  assign n1528_o = x == 9'b101101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:402:13  */
  assign n1531_o = x == 9'b101101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:403:13  */
  assign n1534_o = x == 9'b101101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:404:13  */
  assign n1537_o = x == 9'b101110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:405:13  */
  assign n1540_o = x == 9'b101110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:406:13  */
  assign n1543_o = x == 9'b101110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:407:13  */
  assign n1546_o = x == 9'b101110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:408:13  */
  assign n1549_o = x == 9'b101110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:409:13  */
  assign n1552_o = x == 9'b101110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:410:13  */
  assign n1555_o = x == 9'b101110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:411:13  */
  assign n1558_o = x == 9'b101110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:412:13  */
  assign n1561_o = x == 9'b101111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:413:13  */
  assign n1564_o = x == 9'b101111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:414:13  */
  assign n1567_o = x == 9'b101111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:415:13  */
  assign n1570_o = x == 9'b101111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:416:13  */
  assign n1573_o = x == 9'b101111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:417:13  */
  assign n1576_o = x == 9'b101111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:418:13  */
  assign n1579_o = x == 9'b101111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:419:13  */
  assign n1582_o = x == 9'b101111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:420:13  */
  assign n1585_o = x == 9'b110000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:421:13  */
  assign n1588_o = x == 9'b110000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:422:13  */
  assign n1591_o = x == 9'b110000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:423:13  */
  assign n1594_o = x == 9'b110000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:424:13  */
  assign n1597_o = x == 9'b110000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:425:13  */
  assign n1600_o = x == 9'b110000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:426:13  */
  assign n1603_o = x == 9'b110000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:427:13  */
  assign n1606_o = x == 9'b110000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:428:13  */
  assign n1609_o = x == 9'b110001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:429:13  */
  assign n1612_o = x == 9'b110001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:430:13  */
  assign n1615_o = x == 9'b110001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:431:13  */
  assign n1618_o = x == 9'b110001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:432:13  */
  assign n1621_o = x == 9'b110001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:433:13  */
  assign n1624_o = x == 9'b110001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:434:13  */
  assign n1627_o = x == 9'b110001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:435:13  */
  assign n1630_o = x == 9'b110001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:436:13  */
  assign n1633_o = x == 9'b110010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:437:13  */
  assign n1636_o = x == 9'b110010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:438:13  */
  assign n1639_o = x == 9'b110010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:439:13  */
  assign n1642_o = x == 9'b110010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:440:13  */
  assign n1645_o = x == 9'b110010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:441:13  */
  assign n1648_o = x == 9'b110010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:442:13  */
  assign n1651_o = x == 9'b110010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:443:13  */
  assign n1654_o = x == 9'b110010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:444:13  */
  assign n1657_o = x == 9'b110011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:445:13  */
  assign n1660_o = x == 9'b110011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:446:13  */
  assign n1663_o = x == 9'b110011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:447:13  */
  assign n1666_o = x == 9'b110011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:448:13  */
  assign n1669_o = x == 9'b110011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:449:13  */
  assign n1672_o = x == 9'b110011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:450:13  */
  assign n1675_o = x == 9'b110011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:451:13  */
  assign n1678_o = x == 9'b110011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:452:13  */
  assign n1681_o = x == 9'b110100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:453:13  */
  assign n1684_o = x == 9'b110100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:454:13  */
  assign n1687_o = x == 9'b110100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:455:13  */
  assign n1690_o = x == 9'b110100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:456:13  */
  assign n1693_o = x == 9'b110100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:457:13  */
  assign n1696_o = x == 9'b110100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:458:13  */
  assign n1699_o = x == 9'b110100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:459:13  */
  assign n1702_o = x == 9'b110100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:460:13  */
  assign n1705_o = x == 9'b110101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:461:13  */
  assign n1708_o = x == 9'b110101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:462:13  */
  assign n1711_o = x == 9'b110101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:463:13  */
  assign n1714_o = x == 9'b110101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:464:13  */
  assign n1717_o = x == 9'b110101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:465:13  */
  assign n1720_o = x == 9'b110101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:466:13  */
  assign n1723_o = x == 9'b110101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:467:13  */
  assign n1726_o = x == 9'b110101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:468:13  */
  assign n1729_o = x == 9'b110110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:469:13  */
  assign n1732_o = x == 9'b110110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:470:13  */
  assign n1735_o = x == 9'b110110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:471:13  */
  assign n1738_o = x == 9'b110110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:472:13  */
  assign n1741_o = x == 9'b110110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:473:13  */
  assign n1744_o = x == 9'b110110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:474:13  */
  assign n1747_o = x == 9'b110110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:475:13  */
  assign n1750_o = x == 9'b110110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:476:13  */
  assign n1753_o = x == 9'b110111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:477:13  */
  assign n1756_o = x == 9'b110111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:478:13  */
  assign n1759_o = x == 9'b110111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:479:13  */
  assign n1762_o = x == 9'b110111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:480:13  */
  assign n1765_o = x == 9'b110111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:481:13  */
  assign n1768_o = x == 9'b110111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:482:13  */
  assign n1771_o = x == 9'b110111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:483:13  */
  assign n1774_o = x == 9'b110111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:484:13  */
  assign n1777_o = x == 9'b111000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:485:13  */
  assign n1780_o = x == 9'b111000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:486:13  */
  assign n1783_o = x == 9'b111000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:487:13  */
  assign n1786_o = x == 9'b111000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:488:13  */
  assign n1789_o = x == 9'b111000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:489:13  */
  assign n1792_o = x == 9'b111000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:490:13  */
  assign n1795_o = x == 9'b111000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:491:13  */
  assign n1798_o = x == 9'b111000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:492:13  */
  assign n1801_o = x == 9'b111001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:493:13  */
  assign n1804_o = x == 9'b111001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:494:13  */
  assign n1807_o = x == 9'b111001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:495:13  */
  assign n1810_o = x == 9'b111001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:496:13  */
  assign n1813_o = x == 9'b111001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:497:13  */
  assign n1816_o = x == 9'b111001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:498:13  */
  assign n1819_o = x == 9'b111001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:499:13  */
  assign n1822_o = x == 9'b111001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:500:13  */
  assign n1825_o = x == 9'b111010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:501:13  */
  assign n1828_o = x == 9'b111010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:502:13  */
  assign n1831_o = x == 9'b111010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:503:13  */
  assign n1834_o = x == 9'b111010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:504:13  */
  assign n1837_o = x == 9'b111010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:505:13  */
  assign n1840_o = x == 9'b111010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:506:13  */
  assign n1843_o = x == 9'b111010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:507:13  */
  assign n1846_o = x == 9'b111010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:508:13  */
  assign n1849_o = x == 9'b111011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:509:13  */
  assign n1852_o = x == 9'b111011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:510:13  */
  assign n1855_o = x == 9'b111011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:511:13  */
  assign n1858_o = x == 9'b111011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:512:13  */
  assign n1861_o = x == 9'b111011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:513:13  */
  assign n1864_o = x == 9'b111011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:514:13  */
  assign n1867_o = x == 9'b111011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:515:13  */
  assign n1870_o = x == 9'b111011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:516:13  */
  assign n1873_o = x == 9'b111100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:517:13  */
  assign n1876_o = x == 9'b111100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:518:13  */
  assign n1879_o = x == 9'b111100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:519:13  */
  assign n1882_o = x == 9'b111100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:520:13  */
  assign n1885_o = x == 9'b111100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:521:13  */
  assign n1888_o = x == 9'b111100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:522:13  */
  assign n1891_o = x == 9'b111100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:523:13  */
  assign n1894_o = x == 9'b111100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:524:13  */
  assign n1897_o = x == 9'b111101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:525:13  */
  assign n1900_o = x == 9'b111101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:526:13  */
  assign n1903_o = x == 9'b111101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:527:13  */
  assign n1906_o = x == 9'b111101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:528:13  */
  assign n1909_o = x == 9'b111101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:529:13  */
  assign n1912_o = x == 9'b111101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:530:13  */
  assign n1915_o = x == 9'b111101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:531:13  */
  assign n1918_o = x == 9'b111101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:532:13  */
  assign n1921_o = x == 9'b111110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:533:13  */
  assign n1924_o = x == 9'b111110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:534:13  */
  assign n1927_o = x == 9'b111110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:535:13  */
  assign n1930_o = x == 9'b111110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:536:13  */
  assign n1933_o = x == 9'b111110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:537:13  */
  assign n1936_o = x == 9'b111110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:538:13  */
  assign n1939_o = x == 9'b111110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:539:13  */
  assign n1942_o = x == 9'b111110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:540:13  */
  assign n1945_o = x == 9'b111111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:541:13  */
  assign n1948_o = x == 9'b111111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:542:13  */
  assign n1951_o = x == 9'b111111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:543:13  */
  assign n1954_o = x == 9'b111111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:544:13  */
  assign n1957_o = x == 9'b111111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:545:13  */
  assign n1960_o = x == 9'b111111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:546:13  */
  assign n1963_o = x == 9'b111111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:547:13  */
  assign n1966_o = x == 9'b111111111;
  assign n1968_o = {n1966_o, n1963_o, n1960_o, n1957_o, n1954_o, n1951_o, n1948_o, n1945_o, n1942_o, n1939_o, n1936_o, n1933_o, n1930_o, n1927_o, n1924_o, n1921_o, n1918_o, n1915_o, n1912_o, n1909_o, n1906_o, n1903_o, n1900_o, n1897_o, n1894_o, n1891_o, n1888_o, n1885_o, n1882_o, n1879_o, n1876_o, n1873_o, n1870_o, n1867_o, n1864_o, n1861_o, n1858_o, n1855_o, n1852_o, n1849_o, n1846_o, n1843_o, n1840_o, n1837_o, n1834_o, n1831_o, n1828_o, n1825_o, n1822_o, n1819_o, n1816_o, n1813_o, n1810_o, n1807_o, n1804_o, n1801_o, n1798_o, n1795_o, n1792_o, n1789_o, n1786_o, n1783_o, n1780_o, n1777_o, n1774_o, n1771_o, n1768_o, n1765_o, n1762_o, n1759_o, n1756_o, n1753_o, n1750_o, n1747_o, n1744_o, n1741_o, n1738_o, n1735_o, n1732_o, n1729_o, n1726_o, n1723_o, n1720_o, n1717_o, n1714_o, n1711_o, n1708_o, n1705_o, n1702_o, n1699_o, n1696_o, n1693_o, n1690_o, n1687_o, n1684_o, n1681_o, n1678_o, n1675_o, n1672_o, n1669_o, n1666_o, n1663_o, n1660_o, n1657_o, n1654_o, n1651_o, n1648_o, n1645_o, n1642_o, n1639_o, n1636_o, n1633_o, n1630_o, n1627_o, n1624_o, n1621_o, n1618_o, n1615_o, n1612_o, n1609_o, n1606_o, n1603_o, n1600_o, n1597_o, n1594_o, n1591_o, n1588_o, n1585_o, n1582_o, n1579_o, n1576_o, n1573_o, n1570_o, n1567_o, n1564_o, n1561_o, n1558_o, n1555_o, n1552_o, n1549_o, n1546_o, n1543_o, n1540_o, n1537_o, n1534_o, n1531_o, n1528_o, n1525_o, n1522_o, n1519_o, n1516_o, n1513_o, n1510_o, n1507_o, n1504_o, n1501_o, n1498_o, n1495_o, n1492_o, n1489_o, n1486_o, n1483_o, n1480_o, n1477_o, n1474_o, n1471_o, n1468_o, n1465_o, n1462_o, n1459_o, n1456_o, n1453_o, n1450_o, n1447_o, n1444_o, n1441_o, n1438_o, n1435_o, n1432_o, n1429_o, n1426_o, n1423_o, n1420_o, n1417_o, n1414_o, n1411_o, n1408_o, n1405_o, n1402_o, n1399_o, n1396_o, n1393_o, n1390_o, n1387_o, n1384_o, n1381_o, n1378_o, n1375_o, n1372_o, n1369_o, n1366_o, n1363_o, n1360_o, n1357_o, n1354_o, n1351_o, n1348_o, n1345_o, n1342_o, n1339_o, n1336_o, n1333_o, n1330_o, n1327_o, n1324_o, n1321_o, n1318_o, n1315_o, n1312_o, n1309_o, n1306_o, n1303_o, n1300_o, n1297_o, n1294_o, n1291_o, n1288_o, n1285_o, n1282_o, n1279_o, n1276_o, n1273_o, n1270_o, n1267_o, n1264_o, n1261_o, n1258_o, n1255_o, n1252_o, n1249_o, n1246_o, n1243_o, n1240_o, n1237_o, n1234_o, n1231_o, n1228_o, n1225_o, n1222_o, n1219_o, n1216_o, n1213_o, n1210_o, n1207_o, n1204_o, n1201_o, n1198_o, n1195_o, n1192_o, n1189_o, n1186_o, n1183_o, n1180_o, n1177_o, n1174_o, n1171_o, n1168_o, n1165_o, n1162_o, n1159_o, n1156_o, n1153_o, n1150_o, n1147_o, n1144_o, n1141_o, n1138_o, n1135_o, n1132_o, n1129_o, n1126_o, n1123_o, n1120_o, n1117_o, n1114_o, n1111_o, n1108_o, n1105_o, n1102_o, n1099_o, n1096_o, n1093_o, n1090_o, n1087_o, n1084_o, n1081_o, n1078_o, n1075_o, n1072_o, n1069_o, n1066_o, n1063_o, n1060_o, n1057_o, n1054_o, n1051_o, n1048_o, n1045_o, n1042_o, n1039_o, n1036_o, n1033_o, n1030_o, n1027_o, n1024_o, n1021_o, n1018_o, n1015_o, n1012_o, n1009_o, n1006_o, n1003_o, n1000_o, n997_o, n994_o, n991_o, n988_o, n985_o, n982_o, n979_o, n976_o, n973_o, n970_o, n967_o, n964_o, n961_o, n958_o, n955_o, n952_o, n949_o, n946_o, n943_o, n940_o, n937_o, n934_o, n931_o, n928_o, n925_o, n922_o, n919_o, n916_o, n913_o, n910_o, n907_o, n904_o, n901_o, n898_o, n895_o, n892_o, n889_o, n886_o, n883_o, n880_o, n877_o, n874_o, n871_o, n868_o, n865_o, n862_o, n859_o, n856_o, n853_o, n850_o, n847_o, n844_o, n841_o, n838_o, n835_o, n832_o, n829_o, n826_o, n823_o, n820_o, n817_o, n814_o, n811_o, n808_o, n805_o, n802_o, n799_o, n796_o, n793_o, n790_o, n787_o, n784_o, n781_o, n778_o, n775_o, n772_o, n769_o, n766_o, n763_o, n760_o, n757_o, n754_o, n751_o, n748_o, n745_o, n742_o, n739_o, n736_o, n733_o, n730_o, n727_o, n724_o, n721_o, n718_o, n715_o, n712_o, n709_o, n706_o, n703_o, n700_o, n697_o, n694_o, n691_o, n688_o, n685_o, n682_o, n679_o, n676_o, n673_o, n670_o, n667_o, n664_o, n661_o, n658_o, n655_o, n652_o, n649_o, n646_o, n643_o, n640_o, n637_o, n634_o, n631_o, n628_o, n625_o, n622_o, n619_o, n616_o, n613_o, n610_o, n607_o, n604_o, n601_o, n598_o, n595_o, n592_o, n589_o, n586_o, n583_o, n580_o, n577_o, n574_o, n571_o, n568_o, n565_o, n562_o, n559_o, n556_o, n553_o, n550_o, n547_o, n544_o, n541_o, n538_o, n535_o, n532_o, n529_o, n526_o, n523_o, n520_o, n517_o, n514_o, n511_o, n508_o, n505_o, n502_o, n499_o, n496_o, n493_o, n490_o, n487_o, n484_o, n481_o, n478_o, n475_o, n472_o, n469_o, n466_o, n463_o, n460_o, n457_o, n454_o, n451_o, n448_o, n445_o, n442_o, n439_o, n436_o, n433_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:35:4  */
  always @*
    case (n1968_o)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n1969_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n1969_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n1969_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n1969_o = 3'b000;
      default: n1969_o = 3'bXXX;
    endcase
endmodule

module fdiv #(parameter ID = 1)
  (input wire clk,
   input wire [16:0] X,
   input wire [16:0] Y,
   output wire [16:0] R);
  wire [7:0] fx;
  wire [7:0] fy;
  wire [8:0] expr0;
  wire [8:0] expr0_d1;
  wire [8:0] expr0_d2;
  wire [8:0] expr0_d3;
  wire [8:0] expr0_d4;
  wire [8:0] expr0_d5;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire [3:0] exnxy;
  wire [1:0] exnr0;
  wire [1:0] exnr0_d1;
  wire [1:0] exnr0_d2;
  wire [1:0] exnr0_d3;
  wire [1:0] exnr0_d4;
  wire [1:0] exnr0_d5;
  wire [7:0] d;
  wire [7:0] d_d1;
  wire [7:0] d_d2;
  wire [7:0] d_d3;
  wire [7:0] d_d4;
  wire [8:0] psx;
  wire [10:0] betaw6;
  wire [8:0] sel6;
  wire [2:0] q6;
  wire [2:0] q6_copy5;
  wire [10:0] absq6d;
  wire [10:0] w5;
  wire [10:0] betaw5;
  wire [10:0] betaw5_d1;
  wire [8:0] sel5;
  wire [2:0] q5;
  wire [2:0] q5_copy6;
  wire [2:0] q5_copy6_d1;
  wire [10:0] absq5d;
  wire [10:0] w4;
  wire [10:0] betaw4;
  wire [10:0] betaw4_d1;
  wire [8:0] sel4;
  wire [2:0] q4;
  wire [2:0] q4_copy7;
  wire [2:0] q4_copy7_d1;
  wire [10:0] absq4d;
  wire [10:0] w3;
  wire [10:0] betaw3;
  wire [10:0] betaw3_d1;
  wire [8:0] sel3;
  wire [2:0] q3;
  wire [2:0] q3_d1;
  wire [2:0] q3_copy8;
  wire [10:0] absq3d;
  wire [10:0] absq3d_d1;
  wire [10:0] w2;
  wire [10:0] betaw2;
  wire [8:0] sel2;
  wire [2:0] q2;
  wire [2:0] q2_copy9;
  wire [10:0] absq2d;
  wire [10:0] w1;
  wire [10:0] betaw1;
  wire [10:0] betaw1_d1;
  wire [8:0] sel1;
  wire [2:0] q1;
  wire [2:0] q1_copy10;
  wire [2:0] q1_copy10_d1;
  wire [10:0] absq1d;
  wire [10:0] w0;
  wire [8:0] wfinal;
  wire qm0;
  wire [1:0] qp6;
  wire [1:0] qp6_d1;
  wire [1:0] qp6_d2;
  wire [1:0] qp6_d3;
  wire [1:0] qp6_d4;
  wire [1:0] qm6;
  wire [1:0] qm6_d1;
  wire [1:0] qm6_d2;
  wire [1:0] qm6_d3;
  wire [1:0] qm6_d4;
  wire [1:0] qp5;
  wire [1:0] qp5_d1;
  wire [1:0] qp5_d2;
  wire [1:0] qp5_d3;
  wire [1:0] qm5;
  wire [1:0] qm5_d1;
  wire [1:0] qm5_d2;
  wire [1:0] qm5_d3;
  wire [1:0] qp4;
  wire [1:0] qp4_d1;
  wire [1:0] qp4_d2;
  wire [1:0] qm4;
  wire [1:0] qm4_d1;
  wire [1:0] qm4_d2;
  wire [1:0] qp3;
  wire [1:0] qp3_d1;
  wire [1:0] qp3_d2;
  wire [1:0] qm3;
  wire [1:0] qm3_d1;
  wire [1:0] qm3_d2;
  wire [1:0] qp2;
  wire [1:0] qp2_d1;
  wire [1:0] qm2;
  wire [1:0] qm2_d1;
  wire [1:0] qp1;
  wire [1:0] qm1;
  wire [11:0] qp;
  wire [11:0] qp_d1;
  wire [11:0] qm;
  wire [11:0] qm_d1;
  wire [11:0] quotient;
  wire [9:0] mr;
  wire [7:0] frnorm;
  wire round;
  wire [8:0] expr1;
  wire [15:0] expfrac;
  wire [15:0] expfracr;
  wire [1:0] exnr;
  wire [1:0] exnrfinal;
  wire [6:0] n59_o;
  wire [7:0] n61_o;
  wire [6:0] n62_o;
  wire [7:0] n64_o;
  wire [6:0] n65_o;
  wire [8:0] n67_o;
  wire [6:0] n68_o;
  wire [8:0] n70_o;
  wire [8:0] n71_o;
  wire n72_o;
  wire n73_o;
  wire n74_o;
  wire [1:0] n75_o;
  wire [1:0] n76_o;
  wire [3:0] n77_o;
  wire n80_o;
  wire n83_o;
  wire n85_o;
  wire n86_o;
  wire n88_o;
  wire n89_o;
  wire n92_o;
  wire n94_o;
  wire n95_o;
  wire n97_o;
  wire n98_o;
  wire [2:0] n100_o;
  reg [1:0] n101_o;
  wire [8:0] n103_o;
  wire [10:0] n105_o;
  wire [5:0] n106_o;
  wire [2:0] n107_o;
  wire [8:0] n108_o;
  wire [2:0] selfunctiontable6_n109;
  wire [2:0] selfunctiontable6_y;
  wire [10:0] n113_o;
  wire n115_o;
  wire n117_o;
  wire n118_o;
  wire [9:0] n120_o;
  wire [10:0] n122_o;
  wire n124_o;
  wire n126_o;
  wire n127_o;
  wire [1:0] n129_o;
  reg [10:0] n130_o;
  wire n131_o;
  wire [10:0] n132_o;
  wire n134_o;
  wire [10:0] n135_o;
  reg [10:0] n136_o;
  wire [8:0] n137_o;
  wire [10:0] n139_o;
  wire [5:0] n140_o;
  wire [2:0] n141_o;
  wire [8:0] n142_o;
  wire [2:0] selfunctiontable5_n143;
  wire [2:0] selfunctiontable5_y;
  wire [10:0] n147_o;
  wire n149_o;
  wire n151_o;
  wire n152_o;
  wire [9:0] n154_o;
  wire [10:0] n156_o;
  wire n158_o;
  wire n160_o;
  wire n161_o;
  wire [1:0] n163_o;
  reg [10:0] n164_o;
  wire n165_o;
  wire [10:0] n166_o;
  wire n168_o;
  wire [10:0] n169_o;
  reg [10:0] n170_o;
  wire [8:0] n171_o;
  wire [10:0] n173_o;
  wire [5:0] n174_o;
  wire [2:0] n175_o;
  wire [8:0] n176_o;
  wire [2:0] selfunctiontable4_n177;
  wire [2:0] selfunctiontable4_y;
  wire [10:0] n181_o;
  wire n183_o;
  wire n185_o;
  wire n186_o;
  wire [9:0] n188_o;
  wire [10:0] n190_o;
  wire n192_o;
  wire n194_o;
  wire n195_o;
  wire [1:0] n197_o;
  reg [10:0] n198_o;
  wire n199_o;
  wire [10:0] n200_o;
  wire n202_o;
  wire [10:0] n203_o;
  reg [10:0] n204_o;
  wire [8:0] n205_o;
  wire [10:0] n207_o;
  wire [5:0] n208_o;
  wire [2:0] n209_o;
  wire [8:0] n210_o;
  wire [2:0] selfunctiontable3_n211;
  wire [2:0] selfunctiontable3_y;
  wire [10:0] n215_o;
  wire n217_o;
  wire n219_o;
  wire n220_o;
  wire [9:0] n222_o;
  wire [10:0] n224_o;
  wire n226_o;
  wire n228_o;
  wire n229_o;
  wire [1:0] n231_o;
  reg [10:0] n232_o;
  wire n233_o;
  wire [10:0] n234_o;
  wire n236_o;
  wire [10:0] n237_o;
  reg [10:0] n238_o;
  wire [8:0] n239_o;
  wire [10:0] n241_o;
  wire [5:0] n242_o;
  wire [2:0] n243_o;
  wire [8:0] n244_o;
  wire [2:0] selfunctiontable2_n245;
  wire [2:0] selfunctiontable2_y;
  wire [10:0] n249_o;
  wire n251_o;
  wire n253_o;
  wire n254_o;
  wire [9:0] n256_o;
  wire [10:0] n258_o;
  wire n260_o;
  wire n262_o;
  wire n263_o;
  wire [1:0] n265_o;
  reg [10:0] n266_o;
  wire n267_o;
  wire [10:0] n268_o;
  wire n270_o;
  wire [10:0] n271_o;
  reg [10:0] n272_o;
  wire [8:0] n273_o;
  wire [10:0] n275_o;
  wire [5:0] n276_o;
  wire [2:0] n277_o;
  wire [8:0] n278_o;
  wire [2:0] selfunctiontable1_n279;
  wire [2:0] selfunctiontable1_y;
  wire [10:0] n283_o;
  wire n285_o;
  wire n287_o;
  wire n288_o;
  wire [9:0] n290_o;
  wire [10:0] n292_o;
  wire n294_o;
  wire n296_o;
  wire n297_o;
  wire [1:0] n299_o;
  reg [10:0] n300_o;
  wire n301_o;
  wire [10:0] n302_o;
  wire n304_o;
  wire [10:0] n305_o;
  reg [10:0] n306_o;
  wire [8:0] n307_o;
  wire n308_o;
  wire [1:0] n309_o;
  wire n310_o;
  wire [1:0] n312_o;
  wire [1:0] n313_o;
  wire n314_o;
  wire [1:0] n316_o;
  wire [1:0] n317_o;
  wire n318_o;
  wire [1:0] n320_o;
  wire [1:0] n321_o;
  wire n322_o;
  wire [1:0] n324_o;
  wire [1:0] n325_o;
  wire n326_o;
  wire [1:0] n328_o;
  wire [1:0] n329_o;
  wire n330_o;
  wire [1:0] n332_o;
  wire [3:0] n333_o;
  wire [5:0] n334_o;
  wire [7:0] n335_o;
  wire [9:0] n336_o;
  wire [11:0] n337_o;
  wire n338_o;
  wire [2:0] n339_o;
  wire [4:0] n340_o;
  wire [6:0] n341_o;
  wire [8:0] n342_o;
  wire [10:0] n343_o;
  wire [11:0] n344_o;
  wire [11:0] n345_o;
  wire [9:0] n346_o;
  wire [7:0] n347_o;
  wire n348_o;
  wire [7:0] n349_o;
  wire [7:0] n350_o;
  wire n351_o;
  wire n352_o;
  wire [8:0] n354_o;
  wire [8:0] n355_o;
  wire [6:0] n356_o;
  wire [15:0] n357_o;
  wire [15:0] n359_o;
  wire [15:0] n360_o;
  wire n362_o;
  wire [1:0] n363_o;
  wire [1:0] n365_o;
  wire n367_o;
  wire [1:0] n368_o;
  wire n371_o;
  reg [1:0] n372_o;
  wire [2:0] n373_o;
  wire [13:0] n374_o;
  wire [16:0] n375_o;
  reg [8:0] n376_q;
  reg [8:0] n377_q;
  reg [8:0] n378_q;
  reg [8:0] n379_q;
  reg [8:0] n380_q;
  reg n381_q;
  reg n382_q;
  reg n383_q;
  reg n384_q;
  reg n385_q;
  reg [1:0] n386_q;
  reg [1:0] n387_q;
  reg [1:0] n388_q;
  reg [1:0] n389_q;
  reg [1:0] n390_q;
  reg [7:0] n391_q;
  reg [7:0] n392_q;
  reg [7:0] n393_q;
  reg [7:0] n394_q;
  reg [10:0] n395_q;
  reg [2:0] n396_q;
  reg [10:0] n397_q;
  reg [2:0] n398_q;
  reg [10:0] n399_q;
  reg [2:0] n400_q;
  reg [10:0] n401_q;
  reg [10:0] n402_q;
  reg [2:0] n403_q;
  reg [1:0] n404_q;
  reg [1:0] n405_q;
  reg [1:0] n406_q;
  reg [1:0] n407_q;
  reg [1:0] n408_q;
  reg [1:0] n409_q;
  reg [1:0] n410_q;
  reg [1:0] n411_q;
  reg [1:0] n412_q;
  reg [1:0] n413_q;
  reg [1:0] n414_q;
  reg [1:0] n415_q;
  reg [1:0] n416_q;
  reg [1:0] n417_q;
  reg [1:0] n418_q;
  reg [1:0] n419_q;
  reg [1:0] n420_q;
  reg [1:0] n421_q;
  reg [1:0] n422_q;
  reg [1:0] n423_q;
  reg [1:0] n424_q;
  reg [1:0] n425_q;
  reg [1:0] n426_q;
  reg [1:0] n427_q;
  reg [11:0] n428_q;
  reg [11:0] n429_q;
  assign R = n375_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:588:8  */
  assign fx = n61_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:589:8  */
  assign fy = n64_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:8  */
  assign expr0 = n71_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:15  */
  assign expr0_d1 = n376_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:25  */
  assign expr0_d2 = n377_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:35  */
  assign expr0_d3 = n378_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:45  */
  assign expr0_d4 = n379_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:590:55  */
  assign expr0_d5 = n380_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:8  */
  assign sr = n74_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:12  */
  assign sr_d1 = n381_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:19  */
  assign sr_d2 = n382_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:26  */
  assign sr_d3 = n383_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:33  */
  assign sr_d4 = n384_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:591:40  */
  assign sr_d5 = n385_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:592:8  */
  assign exnxy = n77_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:8  */
  assign exnr0 = n101_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:15  */
  assign exnr0_d1 = n386_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:25  */
  assign exnr0_d2 = n387_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:35  */
  assign exnr0_d3 = n388_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:45  */
  assign exnr0_d4 = n389_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:593:55  */
  assign exnr0_d5 = n390_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:594:8  */
  assign d = fy; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:594:11  */
  assign d_d1 = n391_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:594:17  */
  assign d_d2 = n392_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:594:23  */
  assign d_d3 = n393_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:594:29  */
  assign d_d4 = n394_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:595:8  */
  assign psx = n103_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:596:8  */
  assign betaw6 = n105_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:597:8  */
  assign sel6 = n108_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:598:8  */
  assign q6 = q6_copy5; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:599:8  */
  assign q6_copy5 = selfunctiontable6_n109; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:600:8  */
  assign absq6d = n130_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:601:8  */
  assign w5 = n136_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:602:8  */
  assign betaw5 = n139_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:602:16  */
  assign betaw5_d1 = n395_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:603:8  */
  assign sel5 = n142_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:604:8  */
  assign q5 = q5_copy6_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:605:8  */
  assign q5_copy6 = selfunctiontable5_n143; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:605:18  */
  assign q5_copy6_d1 = n396_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:606:8  */
  assign absq5d = n164_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:607:8  */
  assign w4 = n170_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:608:8  */
  assign betaw4 = n173_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:608:16  */
  assign betaw4_d1 = n397_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:609:8  */
  assign sel4 = n176_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:610:8  */
  assign q4 = q4_copy7_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:611:8  */
  assign q4_copy7 = selfunctiontable4_n177; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:611:18  */
  assign q4_copy7_d1 = n398_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:612:8  */
  assign absq4d = n198_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:613:8  */
  assign w3 = n204_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:614:8  */
  assign betaw3 = n207_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:614:16  */
  assign betaw3_d1 = n399_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:615:8  */
  assign sel3 = n210_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:616:8  */
  assign q3 = q3_copy8; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:616:12  */
  assign q3_d1 = n400_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:617:8  */
  assign q3_copy8 = selfunctiontable3_n211; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:618:8  */
  assign absq3d = n232_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:618:16  */
  assign absq3d_d1 = n401_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:619:8  */
  assign w2 = n238_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:620:8  */
  assign betaw2 = n241_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:621:8  */
  assign sel2 = n244_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:622:8  */
  assign q2 = q2_copy9; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:623:8  */
  assign q2_copy9 = selfunctiontable2_n245; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:624:8  */
  assign absq2d = n266_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:625:8  */
  assign w1 = n272_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:626:8  */
  assign betaw1 = n275_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:626:16  */
  assign betaw1_d1 = n402_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:627:8  */
  assign sel1 = n278_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:628:8  */
  assign q1 = q1_copy10_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:629:8  */
  assign q1_copy10 = selfunctiontable1_n279; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:629:19  */
  assign q1_copy10_d1 = n403_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:630:8  */
  assign absq1d = n300_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:631:8  */
  assign w0 = n306_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:632:8  */
  assign wfinal = n307_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:633:8  */
  assign qm0 = n308_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:634:8  */
  assign qp6 = n309_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:634:13  */
  assign qp6_d1 = n404_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:634:21  */
  assign qp6_d2 = n405_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:634:29  */
  assign qp6_d3 = n406_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:634:37  */
  assign qp6_d4 = n407_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:635:8  */
  assign qm6 = n312_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:635:13  */
  assign qm6_d1 = n408_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:635:21  */
  assign qm6_d2 = n409_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:635:29  */
  assign qm6_d3 = n410_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:635:37  */
  assign qm6_d4 = n411_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:636:8  */
  assign qp5 = n313_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:636:13  */
  assign qp5_d1 = n412_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:636:21  */
  assign qp5_d2 = n413_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:636:29  */
  assign qp5_d3 = n414_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:637:8  */
  assign qm5 = n316_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:637:13  */
  assign qm5_d1 = n415_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:637:21  */
  assign qm5_d2 = n416_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:637:29  */
  assign qm5_d3 = n417_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:638:8  */
  assign qp4 = n317_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:638:13  */
  assign qp4_d1 = n418_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:638:21  */
  assign qp4_d2 = n419_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:639:8  */
  assign qm4 = n320_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:639:13  */
  assign qm4_d1 = n420_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:639:21  */
  assign qm4_d2 = n421_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:640:8  */
  assign qp3 = n321_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:640:13  */
  assign qp3_d1 = n422_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:640:21  */
  assign qp3_d2 = n423_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:641:8  */
  assign qm3 = n324_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:641:13  */
  assign qm3_d1 = n424_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:641:21  */
  assign qm3_d2 = n425_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:642:8  */
  assign qp2 = n325_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:642:13  */
  assign qp2_d1 = n426_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:643:8  */
  assign qm2 = n328_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:643:13  */
  assign qm2_d1 = n427_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:644:8  */
  assign qp1 = n329_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:645:8  */
  assign qm1 = n332_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:646:8  */
  assign qp = n337_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:646:12  */
  assign qp_d1 = n428_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:647:8  */
  assign qm = n344_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:647:12  */
  assign qm_d1 = n429_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:648:8  */
  assign quotient = n345_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:649:8  */
  assign mr = n346_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:650:8  */
  assign frnorm = n349_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:651:8  */
  assign round = n351_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:652:8  */
  assign expr1 = n355_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:653:8  */
  assign expfrac = n357_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:654:8  */
  assign expfracr = n360_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:655:8  */
  assign exnr = n363_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:656:8  */
  assign exnrfinal = n372_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:717:17  */
  assign n59_o = X[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:717:14  */
  assign n61_o = {1'b1, n59_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:718:17  */
  assign n62_o = Y[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:718:14  */
  assign n64_o = {1'b1, n62_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:720:22  */
  assign n65_o = X[13:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:720:19  */
  assign n67_o = {2'b00, n65_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:720:48  */
  assign n68_o = Y[13:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:720:45  */
  assign n70_o = {2'b00, n68_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:720:37  */
  assign n71_o = n67_o - n70_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:721:11  */
  assign n72_o = X[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:721:21  */
  assign n73_o = Y[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:721:16  */
  assign n74_o = n72_o ^ n73_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:723:14  */
  assign n75_o = X[16:15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:723:32  */
  assign n76_o = Y[16:15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:723:29  */
  assign n77_o = {n75_o, n76_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:726:18  */
  assign n80_o = exnxy == 4'b0101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:727:18  */
  assign n83_o = exnxy == 4'b0001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:727:30  */
  assign n85_o = exnxy == 4'b0010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:727:30  */
  assign n86_o = n83_o | n85_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:727:39  */
  assign n88_o = exnxy == 4'b0110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:727:39  */
  assign n89_o = n86_o | n88_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:728:18  */
  assign n92_o = exnxy == 4'b0100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:728:30  */
  assign n94_o = exnxy == 4'b1000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:728:30  */
  assign n95_o = n92_o | n94_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:728:39  */
  assign n97_o = exnxy == 4'b1001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:728:39  */
  assign n98_o = n95_o | n97_o;
  assign n100_o = {n98_o, n89_o, n80_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:724:4  */
  always @*
    case (n100_o)
      3'b100: n101_o = 2'b10;
      3'b010: n101_o = 2'b00;
      3'b001: n101_o = 2'b01;
      default: n101_o = 2'b11;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:731:15  */
  assign n103_o = {1'b0, fx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:732:20  */
  assign n105_o = {2'b00, psx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:733:18  */
  assign n106_o = betaw6[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:733:35  */
  assign n107_o = d[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:733:32  */
  assign n108_o = {n106_o, n107_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:736:23  */
  assign selfunctiontable6_n109 = selfunctiontable6_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:734:4  */
  selfunction_f300_uid4 selfunctiontable6 (
    .x(sel6),
    .y(selfunctiontable6_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:741:16  */
  assign n113_o = {3'b000, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:741:66  */
  assign n115_o = q6 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:741:77  */
  assign n117_o = q6 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:741:77  */
  assign n118_o = n115_o | n117_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:742:15  */
  assign n120_o = {2'b00, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:742:19  */
  assign n122_o = {n120_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:742:52  */
  assign n124_o = q6 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:742:63  */
  assign n126_o = q6 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:742:63  */
  assign n127_o = n124_o | n126_o;
  assign n129_o = {n127_o, n118_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:739:4  */
  always @*
    case (n129_o)
      2'b10: n130_o = n122_o;
      2'b01: n130_o = n113_o;
      default: n130_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:745:11  */
  assign n131_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:746:16  */
  assign n132_o = betaw6 - absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:746:25  */
  assign n134_o = n131_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:747:17  */
  assign n135_o = betaw6 + absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:745:4  */
  always @*
    case (n134_o)
      1'b1: n136_o = n132_o;
      default: n136_o = n135_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:749:16  */
  assign n137_o = w5[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:749:29  */
  assign n139_o = {n137_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:750:18  */
  assign n140_o = betaw5[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:750:35  */
  assign n141_o = d[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:750:32  */
  assign n142_o = {n140_o, n141_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:753:23  */
  assign selfunctiontable5_n143 = selfunctiontable5_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:751:4  */
  selfunction_f300_uid4 selfunctiontable5 (
    .x(sel5),
    .y(selfunctiontable5_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:758:16  */
  assign n147_o = {3'b000, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:758:66  */
  assign n149_o = q5 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:758:77  */
  assign n151_o = q5 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:758:77  */
  assign n152_o = n149_o | n151_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:759:15  */
  assign n154_o = {2'b00, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:759:22  */
  assign n156_o = {n154_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:759:52  */
  assign n158_o = q5 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:759:63  */
  assign n160_o = q5 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:759:63  */
  assign n161_o = n158_o | n160_o;
  assign n163_o = {n161_o, n152_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:756:4  */
  always @*
    case (n163_o)
      2'b10: n164_o = n156_o;
      2'b01: n164_o = n147_o;
      default: n164_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:762:11  */
  assign n165_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:763:19  */
  assign n166_o = betaw5_d1 - absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:763:28  */
  assign n168_o = n165_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:764:20  */
  assign n169_o = betaw5_d1 + absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:762:4  */
  always @*
    case (n168_o)
      1'b1: n170_o = n166_o;
      default: n170_o = n169_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:766:16  */
  assign n171_o = w4[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:766:29  */
  assign n173_o = {n171_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:767:18  */
  assign n174_o = betaw4[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:767:38  */
  assign n175_o = d_d1[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:767:32  */
  assign n176_o = {n174_o, n175_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:770:23  */
  assign selfunctiontable4_n177 = selfunctiontable4_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:768:4  */
  selfunction_f300_uid4 selfunctiontable4 (
    .x(sel4),
    .y(selfunctiontable4_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:775:16  */
  assign n181_o = {3'b000, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:775:66  */
  assign n183_o = q4 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:775:77  */
  assign n185_o = q4 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:775:77  */
  assign n186_o = n183_o | n185_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:776:15  */
  assign n188_o = {2'b00, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:776:22  */
  assign n190_o = {n188_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:776:52  */
  assign n192_o = q4 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:776:63  */
  assign n194_o = q4 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:776:63  */
  assign n195_o = n192_o | n194_o;
  assign n197_o = {n195_o, n186_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:773:4  */
  always @*
    case (n197_o)
      2'b10: n198_o = n190_o;
      2'b01: n198_o = n181_o;
      default: n198_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:779:11  */
  assign n199_o = q4[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:780:19  */
  assign n200_o = betaw4_d1 - absq4d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:780:28  */
  assign n202_o = n199_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:781:20  */
  assign n203_o = betaw4_d1 + absq4d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:779:4  */
  always @*
    case (n202_o)
      1'b1: n204_o = n200_o;
      default: n204_o = n203_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:783:16  */
  assign n205_o = w3[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:783:29  */
  assign n207_o = {n205_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:784:18  */
  assign n208_o = betaw3[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:784:38  */
  assign n209_o = d_d2[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:784:32  */
  assign n210_o = {n208_o, n209_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:787:23  */
  assign selfunctiontable3_n211 = selfunctiontable3_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:785:4  */
  selfunction_f300_uid4 selfunctiontable3 (
    .x(sel3),
    .y(selfunctiontable3_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:792:16  */
  assign n215_o = {3'b000, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:792:66  */
  assign n217_o = q3 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:792:77  */
  assign n219_o = q3 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:792:77  */
  assign n220_o = n217_o | n219_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:793:15  */
  assign n222_o = {2'b00, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:793:22  */
  assign n224_o = {n222_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:793:52  */
  assign n226_o = q3 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:793:63  */
  assign n228_o = q3 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:793:63  */
  assign n229_o = n226_o | n228_o;
  assign n231_o = {n229_o, n220_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:790:4  */
  always @*
    case (n231_o)
      2'b10: n232_o = n224_o;
      2'b01: n232_o = n215_o;
      default: n232_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:796:14  */
  assign n233_o = q3_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:797:19  */
  assign n234_o = betaw3_d1 - absq3d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:797:31  */
  assign n236_o = n233_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:798:20  */
  assign n237_o = betaw3_d1 + absq3d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:796:4  */
  always @*
    case (n236_o)
      1'b1: n238_o = n234_o;
      default: n238_o = n237_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:800:16  */
  assign n239_o = w2[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:800:29  */
  assign n241_o = {n239_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:801:18  */
  assign n242_o = betaw2[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:801:38  */
  assign n243_o = d_d3[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:801:32  */
  assign n244_o = {n242_o, n243_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:804:23  */
  assign selfunctiontable2_n245 = selfunctiontable2_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:802:4  */
  selfunction_f300_uid4 selfunctiontable2 (
    .x(sel2),
    .y(selfunctiontable2_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:809:16  */
  assign n249_o = {3'b000, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:809:66  */
  assign n251_o = q2 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:809:77  */
  assign n253_o = q2 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:809:77  */
  assign n254_o = n251_o | n253_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:810:15  */
  assign n256_o = {2'b00, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:810:22  */
  assign n258_o = {n256_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:810:52  */
  assign n260_o = q2 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:810:63  */
  assign n262_o = q2 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:810:63  */
  assign n263_o = n260_o | n262_o;
  assign n265_o = {n263_o, n254_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:807:4  */
  always @*
    case (n265_o)
      2'b10: n266_o = n258_o;
      2'b01: n266_o = n249_o;
      default: n266_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:813:11  */
  assign n267_o = q2[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:814:16  */
  assign n268_o = betaw2 - absq2d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:814:25  */
  assign n270_o = n267_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:815:17  */
  assign n271_o = betaw2 + absq2d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:813:4  */
  always @*
    case (n270_o)
      1'b1: n272_o = n268_o;
      default: n272_o = n271_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:817:16  */
  assign n273_o = w1[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:817:29  */
  assign n275_o = {n273_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:818:18  */
  assign n276_o = betaw1[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:818:38  */
  assign n277_o = d_d3[6:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:818:32  */
  assign n278_o = {n276_o, n277_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:821:23  */
  assign selfunctiontable1_n279 = selfunctiontable1_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:819:4  */
  selfunction_f300_uid4 selfunctiontable1 (
    .x(sel1),
    .y(selfunctiontable1_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:826:16  */
  assign n283_o = {3'b000, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:826:66  */
  assign n285_o = q1 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:826:77  */
  assign n287_o = q1 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:826:77  */
  assign n288_o = n285_o | n287_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:827:15  */
  assign n290_o = {2'b00, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:827:22  */
  assign n292_o = {n290_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:827:52  */
  assign n294_o = q1 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:827:63  */
  assign n296_o = q1 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:827:63  */
  assign n297_o = n294_o | n296_o;
  assign n299_o = {n297_o, n288_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:824:4  */
  always @*
    case (n299_o)
      2'b10: n300_o = n292_o;
      2'b01: n300_o = n283_o;
      default: n300_o = 11'b00000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:830:11  */
  assign n301_o = q1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:831:19  */
  assign n302_o = betaw1_d1 - absq1d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:831:28  */
  assign n304_o = n301_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:832:20  */
  assign n305_o = betaw1_d1 + absq1d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:830:4  */
  always @*
    case (n304_o)
      1'b1: n306_o = n302_o;
      default: n306_o = n305_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:834:16  */
  assign n307_o = w0[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:835:17  */
  assign n308_o = wfinal[8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:836:18  */
  assign n309_o = q6[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:837:18  */
  assign n310_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:837:22  */
  assign n312_o = {n310_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:838:18  */
  assign n313_o = q5[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:839:18  */
  assign n314_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:839:22  */
  assign n316_o = {n314_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:840:18  */
  assign n317_o = q4[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:841:18  */
  assign n318_o = q4[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:841:22  */
  assign n320_o = {n318_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:842:18  */
  assign n321_o = q3[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:843:18  */
  assign n322_o = q3[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:843:22  */
  assign n324_o = {n322_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:844:18  */
  assign n325_o = q2[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:845:18  */
  assign n326_o = q2[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:845:22  */
  assign n328_o = {n326_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:846:18  */
  assign n329_o = q1[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:847:18  */
  assign n330_o = q1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:847:22  */
  assign n332_o = {n330_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:848:17  */
  assign n333_o = {qp6_d4, qp5_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:848:26  */
  assign n334_o = {n333_o, qp4_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:848:35  */
  assign n335_o = {n334_o, qp3_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:848:44  */
  assign n336_o = {n335_o, qp2_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:848:53  */
  assign n337_o = {n336_o, qp1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:16  */
  assign n338_o = qm6_d4[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:20  */
  assign n339_o = {n338_o, qm5_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:29  */
  assign n340_o = {n339_o, qm4_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:38  */
  assign n341_o = {n340_o, qm3_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:47  */
  assign n342_o = {n341_o, qm2_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:56  */
  assign n343_o = {n342_o, qm1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:849:62  */
  assign n344_o = {n343_o, qm0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:850:22  */
  assign n345_o = qp_d1 - qm_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:854:18  */
  assign n346_o = quotient[10:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:856:19  */
  assign n347_o = mr[8:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:856:40  */
  assign n348_o = mr[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:856:33  */
  assign n349_o = n348_o ? n347_o : n350_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:857:19  */
  assign n350_o = mr[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:858:19  */
  assign n351_o = frnorm[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:859:57  */
  assign n352_o = mr[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:859:53  */
  assign n354_o = {8'b00011111, n352_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:859:22  */
  assign n355_o = expr0_d5 + n354_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:861:29  */
  assign n356_o = frnorm[7:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:861:21  */
  assign n357_o = {expr1, n356_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:862:48  */
  assign n359_o = {15'b000000000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:862:24  */
  assign n360_o = expfrac + n359_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:863:36  */
  assign n362_o = expfracr[15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:863:23  */
  assign n363_o = n362_o ? 2'b00 : n368_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:864:37  */
  assign n365_o = expfracr[15:14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:864:52  */
  assign n367_o = n365_o == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:864:12  */
  assign n368_o = n367_o ? 2'b10 : 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:868:17  */
  assign n371_o = exnr0_d5 == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:866:4  */
  always @*
    case (n371_o)
      1'b1: n372_o = exnr;
      default: n372_o = exnr0_d5;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:870:19  */
  assign n373_o = {exnrfinal, sr_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:870:37  */
  assign n374_o = expfracr[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:870:27  */
  assign n375_o = {n373_o, n374_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n376_q <= expr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n377_q <= expr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n378_q <= expr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n379_q <= expr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n380_q <= expr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n381_q <= sr;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n382_q <= sr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n383_q <= sr_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n384_q <= sr_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n385_q <= sr_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n386_q <= exnr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n387_q <= exnr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n388_q <= exnr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n389_q <= exnr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n390_q <= exnr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n391_q <= d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n392_q <= d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n393_q <= d_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n394_q <= d_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n395_q <= betaw5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n396_q <= q5_copy6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n397_q <= betaw4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n398_q <= q4_copy7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n399_q <= betaw3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n400_q <= q3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n401_q <= absq3d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n402_q <= betaw1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n403_q <= q1_copy10;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n404_q <= qp6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n405_q <= qp6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n406_q <= qp6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n407_q <= qp6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n408_q <= qm6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n409_q <= qm6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n410_q <= qm6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n411_q <= qm6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n412_q <= qp5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n413_q <= qp5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n414_q <= qp5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n415_q <= qm5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n416_q <= qm5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n417_q <= qm5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n418_q <= qp4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n419_q <= qp4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n420_q <= qm4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n421_q <= qm4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n422_q <= qp3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n423_q <= qp3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n424_q <= qm3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n425_q <= qm3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n426_q <= qp2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n427_q <= qm2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n428_q <= qp;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_7_7.vhdl:660:10  */
  always @(posedge clk)
    n429_q <= qm;
endmodule

