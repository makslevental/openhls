module fsqrt#(parameter ID=1)
  (input  clk,
   input  [14:0] X,
   output [14:0] R);
  wire [5:0] fracx;
  wire [5:0] ern0;
  wire [2:0] xsx;
  wire [5:0] ern1;
  wire [5:0] ern1_d1;
  wire [5:0] ern1_d2;
  wire [9:0] fracxnorm;
  wire [1:0] s0;
  wire [9:0] t1;
  wire d1;
  wire [10:0] t1s;
  wire [5:0] t1s_h;
  wire [4:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [9:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [10:0] t2s;
  wire [6:0] t2s_h;
  wire [3:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [9:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [10:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [2:0] t3s_l;
  wire [2:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [9:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [10:0] t4s;
  wire [8:0] t4s_h;
  wire [1:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [9:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [10:0] t5s;
  wire [9:0] t5s_h;
  wire t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [9:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [10:0] t6s;
  wire [10:0] t6s_h;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [9:0] t7;
  wire [7:0] s6;
  wire d8;
  wire [8:0] mr;
  wire [5:0] fr;
  wire [5:0] fr_d1;
  wire round;
  wire round_d1;
  wire [5:0] frrnd;
  wire [11:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [5:0] n16_o;
  wire [4:0] n17_o;
  wire [5:0] n19_o;
  wire [2:0] n20_o;
  wire [5:0] n22_o;
  wire n23_o;
  wire [5:0] n24_o;
  wire [5:0] n25_o;
  wire [6:0] n27_o;
  wire [9:0] n29_o;
  wire n30_o;
  wire n31_o;
  wire [9:0] n32_o;
  wire [7:0] n34_o;
  wire [9:0] n36_o;
  wire [3:0] n38_o;
  wire [3:0] n40_o;
  wire [5:0] n41_o;
  wire [9:0] n42_o;
  wire n43_o;
  wire n44_o;
  wire [10:0] n46_o;
  wire [5:0] n47_o;
  wire [4:0] n48_o;
  wire [2:0] n50_o;
  wire [3:0] n51_o;
  wire n52_o;
  wire [4:0] n53_o;
  wire [5:0] n55_o;
  wire [5:0] n56_o;
  wire [5:0] n57_o;
  wire [5:0] n58_o;
  wire [4:0] n59_o;
  wire [9:0] n60_o;
  wire [2:0] n61_o;
  wire n62_o;
  wire n63_o;
  wire [10:0] n65_o;
  wire [6:0] n66_o;
  wire [3:0] n67_o;
  wire [3:0] n69_o;
  wire [4:0] n70_o;
  wire n71_o;
  wire [5:0] n72_o;
  wire [6:0] n74_o;
  wire [6:0] n75_o;
  wire [6:0] n76_o;
  wire [6:0] n77_o;
  wire [5:0] n78_o;
  wire [9:0] n79_o;
  wire [3:0] n80_o;
  wire n81_o;
  wire n82_o;
  wire [10:0] n84_o;
  wire [7:0] n85_o;
  wire [2:0] n86_o;
  wire [4:0] n88_o;
  wire [5:0] n89_o;
  wire n90_o;
  wire [6:0] n91_o;
  wire [7:0] n93_o;
  wire [7:0] n94_o;
  wire [7:0] n95_o;
  wire [7:0] n96_o;
  wire [6:0] n97_o;
  wire [9:0] n98_o;
  wire [4:0] n99_o;
  wire n100_o;
  wire n101_o;
  wire [10:0] n103_o;
  wire [8:0] n104_o;
  wire [1:0] n105_o;
  wire [5:0] n107_o;
  wire [6:0] n108_o;
  wire n109_o;
  wire [7:0] n110_o;
  wire [8:0] n112_o;
  wire [8:0] n113_o;
  wire [8:0] n114_o;
  wire [8:0] n115_o;
  wire [7:0] n116_o;
  wire [9:0] n117_o;
  wire [5:0] n118_o;
  wire n119_o;
  wire n120_o;
  wire [10:0] n122_o;
  wire [9:0] n123_o;
  wire n124_o;
  wire [6:0] n126_o;
  wire [7:0] n127_o;
  wire n128_o;
  wire [8:0] n129_o;
  wire [9:0] n131_o;
  wire [9:0] n132_o;
  wire [9:0] n133_o;
  wire [9:0] n134_o;
  wire [8:0] n135_o;
  wire [9:0] n136_o;
  wire [6:0] n137_o;
  wire n138_o;
  wire n139_o;
  wire [10:0] n141_o;
  wire [7:0] n143_o;
  wire [8:0] n144_o;
  wire n145_o;
  wire [9:0] n146_o;
  wire [10:0] n148_o;
  wire [10:0] n149_o;
  wire [10:0] n150_o;
  wire [10:0] n151_o;
  wire [9:0] n152_o;
  wire [7:0] n153_o;
  wire n154_o;
  wire n155_o;
  wire [8:0] n156_o;
  wire [5:0] n157_o;
  wire n158_o;
  wire [5:0] n160_o;
  wire [5:0] n161_o;
  wire [11:0] n162_o;
  wire n165_o;
  wire n168_o;
  wire n171_o;
  wire n174_o;
  wire [3:0] n176_o;
  reg [2:0] n177_o;
  wire [14:0] n178_o;
  reg [5:0] n179_q;
  reg [5:0] n180_q;
  reg n181_q;
  reg [7:0] n182_q;
  reg [2:0] n183_q;
  reg [7:0] n184_q;
  reg [4:0] n185_q;
  reg [5:0] n186_q;
  reg n187_q;
  reg [2:0] n188_q;
  reg [2:0] n189_q;
  assign R = n178_o;
  assign fracx = n16_o; // (signal)
  assign ern0 = n19_o; // (signal)
  assign xsx = n20_o; // (signal)
  assign ern1 = n25_o; // (signal)
  assign ern1_d1 = n179_q; // (signal)
  assign ern1_d2 = n180_q; // (signal)
  assign fracxnorm = n32_o; // (signal)
  assign s0 = 2'b01; // (signal)
  assign t1 = n42_o; // (signal)
  assign d1 = n44_o; // (signal)
  assign t1s = n46_o; // (signal)
  assign t1s_h = n47_o; // (signal)
  assign t1s_l = n48_o; // (signal)
  assign u1 = n55_o; // (signal)
  assign t3_h = n57_o; // (signal)
  assign t2 = n60_o; // (signal)
  assign s1 = n61_o; // (signal)
  assign d2 = n63_o; // (signal)
  assign t2s = n65_o; // (signal)
  assign t2s_h = n66_o; // (signal)
  assign t2s_l = n67_o; // (signal)
  assign u2 = n74_o; // (signal)
  assign t4_h = n76_o; // (signal)
  assign t3 = n79_o; // (signal)
  assign s2 = n80_o; // (signal)
  assign d3 = n82_o; // (signal)
  assign d3_d1 = n181_q; // (signal)
  assign t3s = n84_o; // (signal)
  assign t3s_h = n85_o; // (signal)
  assign t3s_h_d1 = n182_q; // (signal)
  assign t3s_l = n86_o; // (signal)
  assign t3s_l_d1 = n183_q; // (signal)
  assign u3 = n93_o; // (signal)
  assign u3_d1 = n184_q; // (signal)
  assign t5_h = n95_o; // (signal)
  assign t4 = n98_o; // (signal)
  assign s3 = n99_o; // (signal)
  assign s3_d1 = n185_q; // (signal)
  assign d4 = n101_o; // (signal)
  assign t4s = n103_o; // (signal)
  assign t4s_h = n104_o; // (signal)
  assign t4s_l = n105_o; // (signal)
  assign u4 = n112_o; // (signal)
  assign t6_h = n114_o; // (signal)
  assign t5 = n117_o; // (signal)
  assign s4 = n118_o; // (signal)
  assign d5 = n120_o; // (signal)
  assign t5s = n122_o; // (signal)
  assign t5s_h = n123_o; // (signal)
  assign t5s_l = n124_o; // (signal)
  assign u5 = n131_o; // (signal)
  assign t7_h = n133_o; // (signal)
  assign t6 = n136_o; // (signal)
  assign s5 = n137_o; // (signal)
  assign d6 = n139_o; // (signal)
  assign t6s = n141_o; // (signal)
  assign t6s_h = t6s; // (signal)
  assign u6 = n148_o; // (signal)
  assign t8_h = n150_o; // (signal)
  assign t7 = n152_o; // (signal)
  assign s6 = n153_o; // (signal)
  assign d8 = n155_o; // (signal)
  assign mr = n156_o; // (signal)
  assign fr = n157_o; // (signal)
  assign fr_d1 = n186_q; // (signal)
  assign round = n158_o; // (signal)
  assign round_d1 = n187_q; // (signal)
  assign frrnd = n161_o; // (signal)
  assign rn2 = n162_o; // (signal)
  assign xsr = n177_o; // (signal)
  assign xsr_d1 = n188_q; // (signal)
  assign xsr_d2 = n189_q; // (signal)
  assign n16_o = X[5:0];
  assign n17_o = X[11:7];
  assign n19_o = {1'b0, n17_o};
  assign n20_o = X[14:12];
  assign n22_o = ern0 + 6'b001111;
  assign n23_o = X[6];
  assign n24_o = {5'b0, n23_o};  //  uext
  assign n25_o = n22_o + n24_o;
  assign n27_o = {1'b1, fracx};
  assign n29_o = {n27_o, 3'b000};
  assign n30_o = X[6];
  assign n31_o = ~n30_o;
  assign n32_o = n31_o ? n29_o : n36_o;
  assign n34_o = {2'b01, fracx};
  assign n36_o = {n34_o, 2'b00};
  assign n38_o = fracxnorm[9:6];
  assign n40_o = 4'b0111 + n38_o;
  assign n41_o = fracxnorm[5:0];
  assign n42_o = {n40_o, n41_o};
  assign n43_o = t1[9];
  assign n44_o = ~n43_o;
  assign n46_o = {t1, 1'b0};
  assign n47_o = t1s[10:5];
  assign n48_o = t1s[4:0];
  assign n50_o = {1'b0, s0};
  assign n51_o = {n50_o, d1};
  assign n52_o = ~d1;
  assign n53_o = {n51_o, n52_o};
  assign n55_o = {n53_o, 1'b1};
  assign n56_o = t1s_h - u1;
  assign n57_o = d1 ? n56_o : n58_o;
  assign n58_o = t1s_h + u1;
  assign n59_o = t3_h[4:0];
  assign n60_o = {n59_o, t1s_l};
  assign n61_o = {s0, d1};
  assign n62_o = t2[9];
  assign n63_o = ~n62_o;
  assign n65_o = {t2, 1'b0};
  assign n66_o = t2s[10:4];
  assign n67_o = t2s[3:0];
  assign n69_o = {1'b0, s1};
  assign n70_o = {n69_o, d2};
  assign n71_o = ~d2;
  assign n72_o = {n70_o, n71_o};
  assign n74_o = {n72_o, 1'b1};
  assign n75_o = t2s_h - u2;
  assign n76_o = d2 ? n75_o : n77_o;
  assign n77_o = t2s_h + u2;
  assign n78_o = t4_h[5:0];
  assign n79_o = {n78_o, t2s_l};
  assign n80_o = {s1, d2};
  assign n81_o = t3[9];
  assign n82_o = ~n81_o;
  assign n84_o = {t3, 1'b0};
  assign n85_o = t3s[10:3];
  assign n86_o = t3s[2:0];
  assign n88_o = {1'b0, s2};
  assign n89_o = {n88_o, d3};
  assign n90_o = ~d3;
  assign n91_o = {n89_o, n90_o};
  assign n93_o = {n91_o, 1'b1};
  assign n94_o = t3s_h_d1 - u3_d1;
  assign n95_o = d3_d1 ? n94_o : n96_o;
  assign n96_o = t3s_h_d1 + u3_d1;
  assign n97_o = t5_h[6:0];
  assign n98_o = {n97_o, t3s_l_d1};
  assign n99_o = {s2, d3};
  assign n100_o = t4[9];
  assign n101_o = ~n100_o;
  assign n103_o = {t4, 1'b0};
  assign n104_o = t4s[10:2];
  assign n105_o = t4s[1:0];
  assign n107_o = {1'b0, s3_d1};
  assign n108_o = {n107_o, d4};
  assign n109_o = ~d4;
  assign n110_o = {n108_o, n109_o};
  assign n112_o = {n110_o, 1'b1};
  assign n113_o = t4s_h - u4;
  assign n114_o = d4 ? n113_o : n115_o;
  assign n115_o = t4s_h + u4;
  assign n116_o = t6_h[7:0];
  assign n117_o = {n116_o, t4s_l};
  assign n118_o = {s3_d1, d4};
  assign n119_o = t5[9];
  assign n120_o = ~n119_o;
  assign n122_o = {t5, 1'b0};
  assign n123_o = t5s[10:1];
  assign n124_o = t5s[0];
  assign n126_o = {1'b0, s4};
  assign n127_o = {n126_o, d5};
  assign n128_o = ~d5;
  assign n129_o = {n127_o, n128_o};
  assign n131_o = {n129_o, 1'b1};
  assign n132_o = t5s_h - u5;
  assign n133_o = d5 ? n132_o : n134_o;
  assign n134_o = t5s_h + u5;
  assign n135_o = t7_h[8:0];
  assign n136_o = {n135_o, t5s_l};
  assign n137_o = {s4, d5};
  assign n138_o = t6[9];
  assign n139_o = ~n138_o;
  assign n141_o = {t6, 1'b0};
  assign n143_o = {1'b0, s5};
  assign n144_o = {n143_o, d6};
  assign n145_o = ~d6;
  assign n146_o = {n144_o, n145_o};
  assign n148_o = {n146_o, 1'b1};
  assign n149_o = t6s_h - u6;
  assign n150_o = d6 ? n149_o : n151_o;
  assign n151_o = t6s_h + u6;
  assign n152_o = t8_h[9:0];
  assign n153_o = {s5, d6};
  assign n154_o = t7[9];
  assign n155_o = ~n154_o;
  assign n156_o = {s6, d8};
  assign n157_o = mr[6:1];
  assign n158_o = mr[0];
  assign n160_o = {5'b00000, round_d1};
  assign n161_o = fr_d1 + n160_o;
  assign n162_o = {ern1_d2, frrnd};
  assign n165_o = xsx == 3'b010;
  assign n168_o = xsx == 3'b100;
  assign n171_o = xsx == 3'b000;
  assign n174_o = xsx == 3'b001;
  assign n176_o = {n174_o, n171_o, n168_o, n165_o};
  always @*
    case (n176_o)
      4'b1000: n177_o = 3'b001;
      4'b0100: n177_o = 3'b000;
      4'b0010: n177_o = 3'b100;
      4'b0001: n177_o = 3'b010;
      default: n177_o = 3'b110;
    endcase
  assign n178_o = {xsr_d2, rn2};
  always @(posedge clk)
    n179_q <= ern1;
  always @(posedge clk)
    n180_q <= ern1_d1;
  always @(posedge clk)
    n181_q <= d3;
  always @(posedge clk)
    n182_q <= t3s_h;
  always @(posedge clk)
    n183_q <= t3s_l;
  always @(posedge clk)
    n184_q <= u3;
  always @(posedge clk)
    n185_q <= s3;
  always @(posedge clk)
    n186_q <= fr;
  always @(posedge clk)
    n187_q <= round;
  always @(posedge clk)
    n188_q <= xsr;
  always @(posedge clk)
    n189_q <= xsr_d1;
endmodule

