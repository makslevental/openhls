module fsqrt#(parameter ID=1)
  (input  clk,
   input  [16:0] X,
   output [16:0] R);
  wire [9:0] fracx;
  wire [3:0] ern0;
  wire [2:0] xsx;
  wire [3:0] ern1;
  wire [3:0] ern1_d1;
  wire [3:0] ern1_d2;
  wire [3:0] ern1_d3;
  wire [13:0] fracxnorm;
  wire [1:0] s0;
  wire [13:0] t1;
  wire d1;
  wire [14:0] t1s;
  wire [5:0] t1s_h;
  wire [8:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [13:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [14:0] t2s;
  wire [6:0] t2s_h;
  wire [7:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [13:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [14:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [6:0] t3s_l;
  wire [6:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [13:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [14:0] t4s;
  wire [8:0] t4s_h;
  wire [5:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [13:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [14:0] t5s;
  wire [9:0] t5s_h;
  wire [4:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [13:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [14:0] t6s;
  wire [10:0] t6s_h;
  wire [3:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [13:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [14:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire [2:0] t7s_l;
  wire [2:0] t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [13:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [14:0] t8s;
  wire [12:0] t8s_h;
  wire [1:0] t8s_l;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [13:0] t9;
  wire [9:0] s8;
  wire d9;
  wire [14:0] t9s;
  wire [13:0] t9s_h;
  wire t9s_l;
  wire [13:0] u9;
  wire [13:0] t11_h;
  wire [13:0] t10;
  wire [10:0] s9;
  wire d10;
  wire d10_d1;
  wire [14:0] t10s;
  wire [14:0] t10s_h;
  wire [14:0] t10s_h_d1;
  wire [14:0] u10;
  wire [14:0] u10_d1;
  wire [14:0] t12_h;
  wire [13:0] t11;
  wire [11:0] s10;
  wire [11:0] s10_d1;
  wire d12;
  wire [12:0] mr;
  wire [9:0] fr;
  wire round;
  wire [9:0] frrnd;
  wire [13:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [2:0] xsr_d3;
  wire [9:0] n25_o;
  wire [2:0] n26_o;
  wire [3:0] n28_o;
  wire [2:0] n29_o;
  wire [3:0] n31_o;
  wire n32_o;
  wire [3:0] n33_o;
  wire [3:0] n34_o;
  wire [10:0] n36_o;
  wire [13:0] n38_o;
  wire n39_o;
  wire n40_o;
  wire [13:0] n41_o;
  wire [11:0] n43_o;
  wire [13:0] n45_o;
  wire [3:0] n47_o;
  wire [3:0] n49_o;
  wire [9:0] n50_o;
  wire [13:0] n51_o;
  wire n52_o;
  wire n53_o;
  wire [14:0] n55_o;
  wire [5:0] n56_o;
  wire [8:0] n57_o;
  wire [2:0] n59_o;
  wire [3:0] n60_o;
  wire n61_o;
  wire [4:0] n62_o;
  wire [5:0] n64_o;
  wire [5:0] n65_o;
  wire [5:0] n66_o;
  wire [5:0] n67_o;
  wire [4:0] n68_o;
  wire [13:0] n69_o;
  wire [2:0] n70_o;
  wire n71_o;
  wire n72_o;
  wire [14:0] n74_o;
  wire [6:0] n75_o;
  wire [7:0] n76_o;
  wire [3:0] n78_o;
  wire [4:0] n79_o;
  wire n80_o;
  wire [5:0] n81_o;
  wire [6:0] n83_o;
  wire [6:0] n84_o;
  wire [6:0] n85_o;
  wire [6:0] n86_o;
  wire [5:0] n87_o;
  wire [13:0] n88_o;
  wire [3:0] n89_o;
  wire n90_o;
  wire n91_o;
  wire [14:0] n93_o;
  wire [7:0] n94_o;
  wire [6:0] n95_o;
  wire [4:0] n97_o;
  wire [5:0] n98_o;
  wire n99_o;
  wire [6:0] n100_o;
  wire [7:0] n102_o;
  wire [7:0] n103_o;
  wire [7:0] n104_o;
  wire [7:0] n105_o;
  wire [6:0] n106_o;
  wire [13:0] n107_o;
  wire [4:0] n108_o;
  wire n109_o;
  wire n110_o;
  wire [14:0] n112_o;
  wire [8:0] n113_o;
  wire [5:0] n114_o;
  wire [5:0] n116_o;
  wire [6:0] n117_o;
  wire n118_o;
  wire [7:0] n119_o;
  wire [8:0] n121_o;
  wire [8:0] n122_o;
  wire [8:0] n123_o;
  wire [8:0] n124_o;
  wire [7:0] n125_o;
  wire [13:0] n126_o;
  wire [5:0] n127_o;
  wire n128_o;
  wire n129_o;
  wire [14:0] n131_o;
  wire [9:0] n132_o;
  wire [4:0] n133_o;
  wire [6:0] n135_o;
  wire [7:0] n136_o;
  wire n137_o;
  wire [8:0] n138_o;
  wire [9:0] n140_o;
  wire [9:0] n141_o;
  wire [9:0] n142_o;
  wire [9:0] n143_o;
  wire [8:0] n144_o;
  wire [13:0] n145_o;
  wire [6:0] n146_o;
  wire n147_o;
  wire n148_o;
  wire [14:0] n150_o;
  wire [10:0] n151_o;
  wire [3:0] n152_o;
  wire [7:0] n154_o;
  wire [8:0] n155_o;
  wire n156_o;
  wire [9:0] n157_o;
  wire [10:0] n159_o;
  wire [10:0] n160_o;
  wire [10:0] n161_o;
  wire [10:0] n162_o;
  wire [9:0] n163_o;
  wire [13:0] n164_o;
  wire [7:0] n165_o;
  wire n166_o;
  wire n167_o;
  wire [14:0] n169_o;
  wire [11:0] n170_o;
  wire [2:0] n171_o;
  wire [8:0] n173_o;
  wire [9:0] n174_o;
  wire n175_o;
  wire [10:0] n176_o;
  wire [11:0] n178_o;
  wire [11:0] n179_o;
  wire [11:0] n180_o;
  wire [11:0] n181_o;
  wire [10:0] n182_o;
  wire [13:0] n183_o;
  wire [8:0] n184_o;
  wire n185_o;
  wire n186_o;
  wire [14:0] n188_o;
  wire [12:0] n189_o;
  wire [1:0] n190_o;
  wire [9:0] n192_o;
  wire [10:0] n193_o;
  wire n194_o;
  wire [11:0] n195_o;
  wire [12:0] n197_o;
  wire [12:0] n198_o;
  wire [12:0] n199_o;
  wire [12:0] n200_o;
  wire [11:0] n201_o;
  wire [13:0] n202_o;
  wire [9:0] n203_o;
  wire n204_o;
  wire n205_o;
  wire [14:0] n207_o;
  wire [13:0] n208_o;
  wire n209_o;
  wire [10:0] n211_o;
  wire [11:0] n212_o;
  wire n213_o;
  wire [12:0] n214_o;
  wire [13:0] n216_o;
  wire [13:0] n217_o;
  wire [13:0] n218_o;
  wire [13:0] n219_o;
  wire [12:0] n220_o;
  wire [13:0] n221_o;
  wire [10:0] n222_o;
  wire n223_o;
  wire n224_o;
  wire [14:0] n226_o;
  wire [11:0] n228_o;
  wire [12:0] n229_o;
  wire n230_o;
  wire [13:0] n231_o;
  wire [14:0] n233_o;
  wire [14:0] n234_o;
  wire [14:0] n235_o;
  wire [14:0] n236_o;
  wire [13:0] n237_o;
  wire [11:0] n238_o;
  wire n239_o;
  wire n240_o;
  wire [12:0] n241_o;
  wire [9:0] n242_o;
  wire n243_o;
  wire [9:0] n245_o;
  wire [9:0] n246_o;
  wire [13:0] n247_o;
  wire n250_o;
  wire n253_o;
  wire n256_o;
  wire n259_o;
  wire [3:0] n261_o;
  reg [2:0] n262_o;
  wire [16:0] n263_o;
  reg [3:0] n264_q;
  reg [3:0] n265_q;
  reg [3:0] n266_q;
  reg n267_q;
  reg [7:0] n268_q;
  reg [6:0] n269_q;
  reg [7:0] n270_q;
  reg [4:0] n271_q;
  reg n272_q;
  reg [11:0] n273_q;
  reg [2:0] n274_q;
  reg [11:0] n275_q;
  reg [8:0] n276_q;
  reg n277_q;
  reg [14:0] n278_q;
  reg [14:0] n279_q;
  reg [11:0] n280_q;
  reg [2:0] n281_q;
  reg [2:0] n282_q;
  reg [2:0] n283_q;
  assign R = n263_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:30:8  */
  assign fracx = n25_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:31:8  */
  assign ern0 = n28_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:32:8  */
  assign xsx = n29_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:33:8  */
  assign ern1 = n34_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:33:14  */
  assign ern1_d1 = n264_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:33:23  */
  assign ern1_d2 = n265_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:33:32  */
  assign ern1_d3 = n266_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:34:8  */
  assign fracxnorm = n41_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:36:8  */
  assign t1 = n51_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:37:8  */
  assign d1 = n53_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:38:8  */
  assign t1s = n55_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:39:8  */
  assign t1s_h = n56_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:40:8  */
  assign t1s_l = n57_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:41:8  */
  assign u1 = n64_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:42:8  */
  assign t3_h = n66_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:43:8  */
  assign t2 = n69_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:44:8  */
  assign s1 = n70_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:45:8  */
  assign d2 = n72_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:46:8  */
  assign t2s = n74_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:47:8  */
  assign t2s_h = n75_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:48:8  */
  assign t2s_l = n76_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:49:8  */
  assign u2 = n83_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:50:8  */
  assign t4_h = n85_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:51:8  */
  assign t3 = n88_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:52:8  */
  assign s2 = n89_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:53:8  */
  assign d3 = n91_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:53:12  */
  assign d3_d1 = n267_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:54:8  */
  assign t3s = n93_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:55:8  */
  assign t3s_h = n94_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:55:15  */
  assign t3s_h_d1 = n268_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:56:8  */
  assign t3s_l = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:56:15  */
  assign t3s_l_d1 = n269_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:57:8  */
  assign u3 = n102_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:57:12  */
  assign u3_d1 = n270_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:58:8  */
  assign t5_h = n104_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:59:8  */
  assign t4 = n107_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:60:8  */
  assign s3 = n108_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:60:12  */
  assign s3_d1 = n271_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:61:8  */
  assign d4 = n110_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:62:8  */
  assign t4s = n112_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:63:8  */
  assign t4s_h = n113_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:64:8  */
  assign t4s_l = n114_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:65:8  */
  assign u4 = n121_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:66:8  */
  assign t6_h = n123_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:67:8  */
  assign t5 = n126_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:68:8  */
  assign s4 = n127_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:69:8  */
  assign d5 = n129_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:70:8  */
  assign t5s = n131_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:71:8  */
  assign t5s_h = n132_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:72:8  */
  assign t5s_l = n133_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:73:8  */
  assign u5 = n140_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:74:8  */
  assign t7_h = n142_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:75:8  */
  assign t6 = n145_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:76:8  */
  assign s5 = n146_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:77:8  */
  assign d6 = n148_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:78:8  */
  assign t6s = n150_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:79:8  */
  assign t6s_h = n151_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:80:8  */
  assign t6s_l = n152_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:81:8  */
  assign u6 = n159_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:82:8  */
  assign t8_h = n161_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:83:8  */
  assign t7 = n164_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:84:8  */
  assign s6 = n165_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:85:8  */
  assign d7 = n167_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:85:12  */
  assign d7_d1 = n272_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:86:8  */
  assign t7s = n169_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:87:8  */
  assign t7s_h = n170_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:87:15  */
  assign t7s_h_d1 = n273_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:88:8  */
  assign t7s_l = n171_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:88:15  */
  assign t7s_l_d1 = n274_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:89:8  */
  assign u7 = n178_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:89:12  */
  assign u7_d1 = n275_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:90:8  */
  assign t9_h = n180_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:91:8  */
  assign t8 = n183_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:92:8  */
  assign s7 = n184_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:92:12  */
  assign s7_d1 = n276_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:93:8  */
  assign d8 = n186_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:94:8  */
  assign t8s = n188_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:95:8  */
  assign t8s_h = n189_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:96:8  */
  assign t8s_l = n190_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:97:8  */
  assign u8 = n197_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:98:8  */
  assign t10_h = n199_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:99:8  */
  assign t9 = n202_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:100:8  */
  assign s8 = n203_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:101:8  */
  assign d9 = n205_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:102:8  */
  assign t9s = n207_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:103:8  */
  assign t9s_h = n208_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:104:8  */
  assign t9s_l = n209_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:105:8  */
  assign u9 = n216_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:106:8  */
  assign t11_h = n218_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:107:8  */
  assign t10 = n221_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:108:8  */
  assign s9 = n222_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:109:8  */
  assign d10 = n224_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:109:13  */
  assign d10_d1 = n277_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:252:18  */
  assign t10s = n226_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:111:8  */
  assign t10s_h = t10s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:111:16  */
  assign t10s_h_d1 = n278_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:112:8  */
  assign u10 = n233_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:112:13  */
  assign u10_d1 = n279_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:113:8  */
  assign t12_h = n235_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:114:8  */
  assign t11 = n237_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:115:8  */
  assign s10 = n238_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:115:13  */
  assign s10_d1 = n280_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:116:8  */
  assign d12 = n240_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:117:8  */
  assign mr = n241_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:118:8  */
  assign fr = n242_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:119:8  */
  assign round = n243_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:120:8  */
  assign frrnd = n246_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:121:8  */
  assign rn2 = n247_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:122:8  */
  assign xsr = n262_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:122:13  */
  assign xsr_d1 = n281_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:122:21  */
  assign xsr_d2 = n282_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:122:29  */
  assign xsr_d3 = n283_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:149:14  */
  assign n25_o = X[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:150:19  */
  assign n26_o = X[13:11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:150:16  */
  assign n28_o = {1'b0, n26_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:151:12  */
  assign n29_o = X[16:14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:152:17  */
  assign n31_o = ern0 + 4'b0011;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:152:51  */
  assign n32_o = X[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:152:48  */
  assign n33_o = {3'b0, n32_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:152:48  */
  assign n34_o = n31_o + n33_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:153:21  */
  assign n36_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:153:29  */
  assign n38_o = {n36_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:153:43  */
  assign n39_o = X[10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:153:48  */
  assign n40_o = ~n39_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:153:37  */
  assign n41_o = n40_o ? n38_o : n45_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:154:15  */
  assign n43_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:154:22  */
  assign n45_o = {n43_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:156:29  */
  assign n47_o = fracxnorm[13:10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:156:18  */
  assign n49_o = 4'b0111 + n47_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:156:56  */
  assign n50_o = fracxnorm[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:156:45  */
  assign n51_o = {n49_o, n50_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:160:16  */
  assign n52_o = t1[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:160:10  */
  assign n53_o = ~n52_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:161:14  */
  assign n55_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:162:16  */
  assign n56_o = t1s[14:9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:163:16  */
  assign n57_o = t1s[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:164:15  */
  assign n59_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:164:20  */
  assign n60_o = {n59_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:164:28  */
  assign n61_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:164:25  */
  assign n62_o = {n60_o, n61_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:164:36  */
  assign n64_o = {n62_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:165:20  */
  assign n65_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:165:25  */
  assign n66_o = d1 ? n65_o : n67_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:166:20  */
  assign n67_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:167:14  */
  assign n68_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:167:27  */
  assign n69_o = {n68_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:168:13  */
  assign n70_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:170:16  */
  assign n71_o = t2[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:170:10  */
  assign n72_o = ~n71_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:171:14  */
  assign n74_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:172:16  */
  assign n75_o = t2s[14:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:173:16  */
  assign n76_o = t2s[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:174:15  */
  assign n78_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:174:20  */
  assign n79_o = {n78_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:174:28  */
  assign n80_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:174:25  */
  assign n81_o = {n79_o, n80_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:174:36  */
  assign n83_o = {n81_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:175:20  */
  assign n84_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:175:25  */
  assign n85_o = d2 ? n84_o : n86_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:176:20  */
  assign n86_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:177:14  */
  assign n87_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:177:27  */
  assign n88_o = {n87_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:178:13  */
  assign n89_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:180:16  */
  assign n90_o = t3[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:180:10  */
  assign n91_o = ~n90_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:181:14  */
  assign n93_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:182:16  */
  assign n94_o = t3s[14:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:183:16  */
  assign n95_o = t3s[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:184:15  */
  assign n97_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:184:20  */
  assign n98_o = {n97_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:184:28  */
  assign n99_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:184:25  */
  assign n100_o = {n98_o, n99_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:184:36  */
  assign n102_o = {n100_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:185:23  */
  assign n103_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:185:31  */
  assign n104_o = d3_d1 ? n103_o : n105_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:186:23  */
  assign n105_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:187:14  */
  assign n106_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:187:27  */
  assign n107_o = {n106_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:188:13  */
  assign n108_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:190:16  */
  assign n109_o = t4[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:190:10  */
  assign n110_o = ~n109_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:191:14  */
  assign n112_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:192:16  */
  assign n113_o = t4s[14:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:193:16  */
  assign n114_o = t4s[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:194:15  */
  assign n116_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:194:23  */
  assign n117_o = {n116_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:194:31  */
  assign n118_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:194:28  */
  assign n119_o = {n117_o, n118_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:194:39  */
  assign n121_o = {n119_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:195:20  */
  assign n122_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:195:25  */
  assign n123_o = d4 ? n122_o : n124_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:196:20  */
  assign n124_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:197:14  */
  assign n125_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:197:27  */
  assign n126_o = {n125_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:198:16  */
  assign n127_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:200:16  */
  assign n128_o = t5[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:200:10  */
  assign n129_o = ~n128_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:201:14  */
  assign n131_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:202:16  */
  assign n132_o = t5s[14:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:203:16  */
  assign n133_o = t5s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:204:15  */
  assign n135_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:204:20  */
  assign n136_o = {n135_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:204:28  */
  assign n137_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:204:25  */
  assign n138_o = {n136_o, n137_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:204:36  */
  assign n140_o = {n138_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:205:20  */
  assign n141_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:205:25  */
  assign n142_o = d5 ? n141_o : n143_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:206:20  */
  assign n143_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:207:14  */
  assign n144_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:207:27  */
  assign n145_o = {n144_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:208:13  */
  assign n146_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:210:16  */
  assign n147_o = t6[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:210:10  */
  assign n148_o = ~n147_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:211:14  */
  assign n150_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:212:16  */
  assign n151_o = t6s[14:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:213:16  */
  assign n152_o = t6s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:214:15  */
  assign n154_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:214:20  */
  assign n155_o = {n154_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:214:28  */
  assign n156_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:214:25  */
  assign n157_o = {n155_o, n156_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:214:36  */
  assign n159_o = {n157_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:215:20  */
  assign n160_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:215:25  */
  assign n161_o = d6 ? n160_o : n162_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:216:20  */
  assign n162_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:217:14  */
  assign n163_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:217:27  */
  assign n164_o = {n163_o, t6s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:218:13  */
  assign n165_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:220:16  */
  assign n166_o = t7[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:220:10  */
  assign n167_o = ~n166_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:221:14  */
  assign n169_o = {t7, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:222:16  */
  assign n170_o = t7s[14:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:223:16  */
  assign n171_o = t7s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:224:15  */
  assign n173_o = {1'b0, s6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:224:20  */
  assign n174_o = {n173_o, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:224:28  */
  assign n175_o = ~d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:224:25  */
  assign n176_o = {n174_o, n175_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:224:36  */
  assign n178_o = {n176_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:225:23  */
  assign n179_o = t7s_h_d1 - u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:225:31  */
  assign n180_o = d7_d1 ? n179_o : n181_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:226:23  */
  assign n181_o = t7s_h_d1 + u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:227:14  */
  assign n182_o = t9_h[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:227:28  */
  assign n183_o = {n182_o, t7s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:228:13  */
  assign n184_o = {s6, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:230:16  */
  assign n185_o = t8[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:230:10  */
  assign n186_o = ~n185_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:231:14  */
  assign n188_o = {t8, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:232:16  */
  assign n189_o = t8s[14:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:233:16  */
  assign n190_o = t8s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:234:15  */
  assign n192_o = {1'b0, s7_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:234:23  */
  assign n193_o = {n192_o, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:234:31  */
  assign n194_o = ~d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:234:28  */
  assign n195_o = {n193_o, n194_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:234:39  */
  assign n197_o = {n195_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:235:21  */
  assign n198_o = t8s_h - u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:235:26  */
  assign n199_o = d8 ? n198_o : n200_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:236:20  */
  assign n200_o = t8s_h + u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:237:15  */
  assign n201_o = t10_h[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:237:29  */
  assign n202_o = {n201_o, t8s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:238:16  */
  assign n203_o = {s7_d1, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:240:16  */
  assign n204_o = t9[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:240:10  */
  assign n205_o = ~n204_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:241:14  */
  assign n207_o = {t9, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:242:16  */
  assign n208_o = t9s[14:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:243:16  */
  assign n209_o = t9s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:244:15  */
  assign n211_o = {1'b0, s8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:244:20  */
  assign n212_o = {n211_o, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:244:28  */
  assign n213_o = ~d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:244:25  */
  assign n214_o = {n212_o, n213_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:244:36  */
  assign n216_o = {n214_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:245:21  */
  assign n217_o = t9s_h - u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:245:26  */
  assign n218_o = d9 ? n217_o : n219_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:246:20  */
  assign n219_o = t9s_h + u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:247:16  */
  assign n220_o = t11_h[12:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:247:30  */
  assign n221_o = {n220_o, t9s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:248:13  */
  assign n222_o = {s8, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:250:18  */
  assign n223_o = t10[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:250:11  */
  assign n224_o = ~n223_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:251:16  */
  assign n226_o = {t10, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:253:16  */
  assign n228_o = {1'b0, s9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:253:21  */
  assign n229_o = {n228_o, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:253:30  */
  assign n230_o = ~d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:253:27  */
  assign n231_o = {n229_o, n230_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:253:39  */
  assign n233_o = {n231_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:254:25  */
  assign n234_o = t10s_h_d1 - u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:254:34  */
  assign n235_o = d10_d1 ? n234_o : n236_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:255:24  */
  assign n236_o = t10s_h_d1 + u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:256:16  */
  assign n237_o = t12_h[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:257:14  */
  assign n238_o = {s9, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:258:18  */
  assign n239_o = t11[13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:258:11  */
  assign n240_o = ~n239_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:259:17  */
  assign n241_o = {s10_d1, d12};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:260:12  */
  assign n242_o = mr[10:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:261:15  */
  assign n243_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:262:39  */
  assign n245_o = {9'b000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:262:16  */
  assign n246_o = fr + n245_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:263:19  */
  assign n247_o = {ern1_d3, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:266:21  */
  assign n250_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:267:21  */
  assign n253_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:268:21  */
  assign n256_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:269:21  */
  assign n259_o = xsx == 3'b001;
  assign n261_o = {n259_o, n256_o, n253_o, n250_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:265:4  */
  always @*
    case (n261_o)
      4'b1000: n262_o = 3'b001;
      4'b0100: n262_o = 3'b000;
      4'b0010: n262_o = 3'b100;
      4'b0001: n262_o = 3'b010;
      default: n262_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:271:16  */
  assign n263_o = {xsr_d3, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n264_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n265_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n266_q <= ern1_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n267_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n268_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n269_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n270_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n271_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n272_q <= d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n273_q <= t7s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n274_q <= t7s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n275_q <= u7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n276_q <= s7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n277_q <= d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n278_q <= t10s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n279_q <= u10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n280_q <= s10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n281_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n282_q <= xsr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_4_10.vhdl:126:10  */
  always @(posedge clk)
    n283_q <= xsr_d2;
endmodule

