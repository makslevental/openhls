module fsqrt#(parameter ID=1)
  (input wire clk,
   input wire [18:0] X,
   output wire [18:0] R);
  wire [10:0] fracx;
  wire [4:0] ern0;
  wire [2:0] xsx;
  wire [4:0] ern1;
  wire [4:0] ern1_d1;
  wire [4:0] ern1_d2;
  wire [4:0] ern1_d3;
  wire [14:0] fracxnorm;
  wire [1:0] s0;
  wire [14:0] t1;
  wire d1;
  wire [15:0] t1s;
  wire [5:0] t1s_h;
  wire [9:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [14:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [15:0] t2s;
  wire [6:0] t2s_h;
  wire [8:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [14:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [15:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [7:0] t3s_l;
  wire [7:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [14:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [15:0] t4s;
  wire [8:0] t4s_h;
  wire [6:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [14:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [15:0] t5s;
  wire [9:0] t5s_h;
  wire [5:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [14:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [15:0] t6s;
  wire [10:0] t6s_h;
  wire [4:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [14:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [15:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire [3:0] t7s_l;
  wire [3:0] t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [14:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [15:0] t8s;
  wire [12:0] t8s_h;
  wire [2:0] t8s_l;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [14:0] t9;
  wire [9:0] s8;
  wire d9;
  wire [15:0] t9s;
  wire [13:0] t9s_h;
  wire [1:0] t9s_l;
  wire [13:0] u9;
  wire [13:0] t11_h;
  wire [14:0] t10;
  wire [10:0] s9;
  wire d10;
  wire d10_d1;
  wire [15:0] t10s;
  wire [14:0] t10s_h;
  wire [14:0] t10s_h_d1;
  wire t10s_l;
  wire t10s_l_d1;
  wire [14:0] u10;
  wire [14:0] u10_d1;
  wire [14:0] t12_h;
  wire [14:0] t11;
  wire [11:0] s10;
  wire [11:0] s10_d1;
  wire d11;
  wire [15:0] t11s;
  wire [15:0] t11s_h;
  wire [15:0] u11;
  wire [15:0] t13_h;
  wire [14:0] t12;
  wire [12:0] s11;
  wire d13;
  wire [13:0] mr;
  wire [10:0] fr;
  wire round;
  wire [10:0] frrnd;
  wire [15:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [2:0] xsr_d3;
  wire [10:0] n26_o;
  wire [3:0] n27_o;
  wire [4:0] n29_o;
  wire [2:0] n30_o;
  wire [4:0] n32_o;
  wire n33_o;
  wire [4:0] n34_o;
  wire [4:0] n35_o;
  wire [11:0] n37_o;
  wire [14:0] n39_o;
  wire n40_o;
  wire n41_o;
  wire [14:0] n42_o;
  wire [12:0] n44_o;
  wire [14:0] n46_o;
  wire [3:0] n48_o;
  wire [3:0] n50_o;
  wire [10:0] n51_o;
  wire [14:0] n52_o;
  wire n53_o;
  wire n54_o;
  wire [15:0] n56_o;
  wire [5:0] n57_o;
  wire [9:0] n58_o;
  wire [2:0] n60_o;
  wire [3:0] n61_o;
  wire n62_o;
  wire [4:0] n63_o;
  wire [5:0] n65_o;
  wire [5:0] n66_o;
  wire [5:0] n67_o;
  wire [5:0] n68_o;
  wire [4:0] n69_o;
  wire [14:0] n70_o;
  wire [2:0] n71_o;
  wire n72_o;
  wire n73_o;
  wire [15:0] n75_o;
  wire [6:0] n76_o;
  wire [8:0] n77_o;
  wire [3:0] n79_o;
  wire [4:0] n80_o;
  wire n81_o;
  wire [5:0] n82_o;
  wire [6:0] n84_o;
  wire [6:0] n85_o;
  wire [6:0] n86_o;
  wire [6:0] n87_o;
  wire [5:0] n88_o;
  wire [14:0] n89_o;
  wire [3:0] n90_o;
  wire n91_o;
  wire n92_o;
  wire [15:0] n94_o;
  wire [7:0] n95_o;
  wire [7:0] n96_o;
  wire [4:0] n98_o;
  wire [5:0] n99_o;
  wire n100_o;
  wire [6:0] n101_o;
  wire [7:0] n103_o;
  wire [7:0] n104_o;
  wire [7:0] n105_o;
  wire [7:0] n106_o;
  wire [6:0] n107_o;
  wire [14:0] n108_o;
  wire [4:0] n109_o;
  wire n110_o;
  wire n111_o;
  wire [15:0] n113_o;
  wire [8:0] n114_o;
  wire [6:0] n115_o;
  wire [5:0] n117_o;
  wire [6:0] n118_o;
  wire n119_o;
  wire [7:0] n120_o;
  wire [8:0] n122_o;
  wire [8:0] n123_o;
  wire [8:0] n124_o;
  wire [8:0] n125_o;
  wire [7:0] n126_o;
  wire [14:0] n127_o;
  wire [5:0] n128_o;
  wire n129_o;
  wire n130_o;
  wire [15:0] n132_o;
  wire [9:0] n133_o;
  wire [5:0] n134_o;
  wire [6:0] n136_o;
  wire [7:0] n137_o;
  wire n138_o;
  wire [8:0] n139_o;
  wire [9:0] n141_o;
  wire [9:0] n142_o;
  wire [9:0] n143_o;
  wire [9:0] n144_o;
  wire [8:0] n145_o;
  wire [14:0] n146_o;
  wire [6:0] n147_o;
  wire n148_o;
  wire n149_o;
  wire [15:0] n151_o;
  wire [10:0] n152_o;
  wire [4:0] n153_o;
  wire [7:0] n155_o;
  wire [8:0] n156_o;
  wire n157_o;
  wire [9:0] n158_o;
  wire [10:0] n160_o;
  wire [10:0] n161_o;
  wire [10:0] n162_o;
  wire [10:0] n163_o;
  wire [9:0] n164_o;
  wire [14:0] n165_o;
  wire [7:0] n166_o;
  wire n167_o;
  wire n168_o;
  wire [15:0] n170_o;
  wire [11:0] n171_o;
  wire [3:0] n172_o;
  wire [8:0] n174_o;
  wire [9:0] n175_o;
  wire n176_o;
  wire [10:0] n177_o;
  wire [11:0] n179_o;
  wire [11:0] n180_o;
  wire [11:0] n181_o;
  wire [11:0] n182_o;
  wire [10:0] n183_o;
  wire [14:0] n184_o;
  wire [8:0] n185_o;
  wire n186_o;
  wire n187_o;
  wire [15:0] n189_o;
  wire [12:0] n190_o;
  wire [2:0] n191_o;
  wire [9:0] n193_o;
  wire [10:0] n194_o;
  wire n195_o;
  wire [11:0] n196_o;
  wire [12:0] n198_o;
  wire [12:0] n199_o;
  wire [12:0] n200_o;
  wire [12:0] n201_o;
  wire [11:0] n202_o;
  wire [14:0] n203_o;
  wire [9:0] n204_o;
  wire n205_o;
  wire n206_o;
  wire [15:0] n208_o;
  wire [13:0] n209_o;
  wire [1:0] n210_o;
  wire [10:0] n212_o;
  wire [11:0] n213_o;
  wire n214_o;
  wire [12:0] n215_o;
  wire [13:0] n217_o;
  wire [13:0] n218_o;
  wire [13:0] n219_o;
  wire [13:0] n220_o;
  wire [12:0] n221_o;
  wire [14:0] n222_o;
  wire [10:0] n223_o;
  wire n224_o;
  wire n225_o;
  wire [15:0] n227_o;
  wire [14:0] n228_o;
  wire n229_o;
  wire [11:0] n231_o;
  wire [12:0] n232_o;
  wire n233_o;
  wire [13:0] n234_o;
  wire [14:0] n236_o;
  wire [14:0] n237_o;
  wire [14:0] n238_o;
  wire [14:0] n239_o;
  wire [13:0] n240_o;
  wire [14:0] n241_o;
  wire [11:0] n242_o;
  wire n243_o;
  wire n244_o;
  wire [15:0] n246_o;
  wire [12:0] n248_o;
  wire [13:0] n249_o;
  wire n250_o;
  wire [14:0] n251_o;
  wire [15:0] n253_o;
  wire [15:0] n254_o;
  wire [15:0] n255_o;
  wire [15:0] n256_o;
  wire [14:0] n257_o;
  wire [12:0] n258_o;
  wire n259_o;
  wire n260_o;
  wire [13:0] n261_o;
  wire [10:0] n262_o;
  wire n263_o;
  wire [10:0] n265_o;
  wire [10:0] n266_o;
  wire [15:0] n267_o;
  wire n270_o;
  wire n273_o;
  wire n276_o;
  wire n279_o;
  wire [3:0] n281_o;
  reg [2:0] n282_o;
  wire [18:0] n283_o;
  reg [4:0] n284_q;
  reg [4:0] n285_q;
  reg [4:0] n286_q;
  reg n287_q;
  reg [7:0] n288_q;
  reg [7:0] n289_q;
  reg [7:0] n290_q;
  reg [4:0] n291_q;
  reg n292_q;
  reg [11:0] n293_q;
  reg [3:0] n294_q;
  reg [11:0] n295_q;
  reg [8:0] n296_q;
  reg n297_q;
  reg [14:0] n298_q;
  reg n299_q;
  reg [14:0] n300_q;
  reg [11:0] n301_q;
  reg [2:0] n302_q;
  reg [2:0] n303_q;
  reg [2:0] n304_q;
  assign R = n283_o;
  assign fracx = n26_o; // (signal)
  assign ern0 = n29_o; // (signal)
  assign xsx = n30_o; // (signal)
  assign ern1 = n35_o; // (signal)
  assign ern1_d1 = n284_q; // (signal)
  assign ern1_d2 = n285_q; // (signal)
  assign ern1_d3 = n286_q; // (signal)
  assign fracxnorm = n42_o; // (signal)
  assign s0 = 2'b01; // (signal)
  assign t1 = n52_o; // (signal)
  assign d1 = n54_o; // (signal)
  assign t1s = n56_o; // (signal)
  assign t1s_h = n57_o; // (signal)
  assign t1s_l = n58_o; // (signal)
  assign u1 = n65_o; // (signal)
  assign t3_h = n67_o; // (signal)
  assign t2 = n70_o; // (signal)
  assign s1 = n71_o; // (signal)
  assign d2 = n73_o; // (signal)
  assign t2s = n75_o; // (signal)
  assign t2s_h = n76_o; // (signal)
  assign t2s_l = n77_o; // (signal)
  assign u2 = n84_o; // (signal)
  assign t4_h = n86_o; // (signal)
  assign t3 = n89_o; // (signal)
  assign s2 = n90_o; // (signal)
  assign d3 = n92_o; // (signal)
  assign d3_d1 = n287_q; // (signal)
  assign t3s = n94_o; // (signal)
  assign t3s_h = n95_o; // (signal)
  assign t3s_h_d1 = n288_q; // (signal)
  assign t3s_l = n96_o; // (signal)
  assign t3s_l_d1 = n289_q; // (signal)
  assign u3 = n103_o; // (signal)
  assign u3_d1 = n290_q; // (signal)
  assign t5_h = n105_o; // (signal)
  assign t4 = n108_o; // (signal)
  assign s3 = n109_o; // (signal)
  assign s3_d1 = n291_q; // (signal)
  assign d4 = n111_o; // (signal)
  assign t4s = n113_o; // (signal)
  assign t4s_h = n114_o; // (signal)
  assign t4s_l = n115_o; // (signal)
  assign u4 = n122_o; // (signal)
  assign t6_h = n124_o; // (signal)
  assign t5 = n127_o; // (signal)
  assign s4 = n128_o; // (signal)
  assign d5 = n130_o; // (signal)
  assign t5s = n132_o; // (signal)
  assign t5s_h = n133_o; // (signal)
  assign t5s_l = n134_o; // (signal)
  assign u5 = n141_o; // (signal)
  assign t7_h = n143_o; // (signal)
  assign t6 = n146_o; // (signal)
  assign s5 = n147_o; // (signal)
  assign d6 = n149_o; // (signal)
  assign t6s = n151_o; // (signal)
  assign t6s_h = n152_o; // (signal)
  assign t6s_l = n153_o; // (signal)
  assign u6 = n160_o; // (signal)
  assign t8_h = n162_o; // (signal)
  assign t7 = n165_o; // (signal)
  assign s6 = n166_o; // (signal)
  assign d7 = n168_o; // (signal)
  assign d7_d1 = n292_q; // (signal)
  assign t7s = n170_o; // (signal)
  assign t7s_h = n171_o; // (signal)
  assign t7s_h_d1 = n293_q; // (signal)
  assign t7s_l = n172_o; // (signal)
  assign t7s_l_d1 = n294_q; // (signal)
  assign u7 = n179_o; // (signal)
  assign u7_d1 = n295_q; // (signal)
  assign t9_h = n181_o; // (signal)
  assign t8 = n184_o; // (signal)
  assign s7 = n185_o; // (signal)
  assign s7_d1 = n296_q; // (signal)
  assign d8 = n187_o; // (signal)
  assign t8s = n189_o; // (signal)
  assign t8s_h = n190_o; // (signal)
  assign t8s_l = n191_o; // (signal)
  assign u8 = n198_o; // (signal)
  assign t10_h = n200_o; // (signal)
  assign t9 = n203_o; // (signal)
  assign s8 = n204_o; // (signal)
  assign d9 = n206_o; // (signal)
  assign t9s = n208_o; // (signal)
  assign t9s_h = n209_o; // (signal)
  assign t9s_l = n210_o; // (signal)
  assign u9 = n217_o; // (signal)
  assign t11_h = n219_o; // (signal)
  assign t10 = n222_o; // (signal)
  assign s9 = n223_o; // (signal)
  assign d10 = n225_o; // (signal)
  assign d10_d1 = n297_q; // (signal)
  assign t10s = n227_o; // (signal)
  assign t10s_h = n228_o; // (signal)
  assign t10s_h_d1 = n298_q; // (signal)
  assign t10s_l = n229_o; // (signal)
  assign t10s_l_d1 = n299_q; // (signal)
  assign u10 = n236_o; // (signal)
  assign u10_d1 = n300_q; // (signal)
  assign t12_h = n238_o; // (signal)
  assign t11 = n241_o; // (signal)
  assign s10 = n242_o; // (signal)
  assign s10_d1 = n301_q; // (signal)
  assign d11 = n244_o; // (signal)
  assign t11s = n246_o; // (signal)
  assign t11s_h = t11s; // (signal)
  assign u11 = n253_o; // (signal)
  assign t13_h = n255_o; // (signal)
  assign t12 = n257_o; // (signal)
  assign s11 = n258_o; // (signal)
  assign d13 = n260_o; // (signal)
  assign mr = n261_o; // (signal)
  assign fr = n262_o; // (signal)
  assign round = n263_o; // (signal)
  assign frrnd = n266_o; // (signal)
  assign rn2 = n267_o; // (signal)
  assign xsr = n282_o; // (signal)
  assign xsr_d1 = n302_q; // (signal)
  assign xsr_d2 = n303_q; // (signal)
  assign xsr_d3 = n304_q; // (signal)
  assign n26_o = X[10:0];
  assign n27_o = X[15:12];
  assign n29_o = {1'b0, n27_o};
  assign n30_o = X[18:16];
  assign n32_o = ern0 + 5'b00111;
  assign n33_o = X[11];
  assign n34_o = {4'b0, n33_o};  //  uext
  assign n35_o = n32_o + n34_o;
  assign n37_o = {1'b1, fracx};
  assign n39_o = {n37_o, 3'b000};
  assign n40_o = X[11];
  assign n41_o = ~n40_o;
  assign n42_o = n41_o ? n39_o : n46_o;
  assign n44_o = {2'b01, fracx};
  assign n46_o = {n44_o, 2'b00};
  assign n48_o = fracxnorm[14:11];
  assign n50_o = 4'b0111 + n48_o;
  assign n51_o = fracxnorm[10:0];
  assign n52_o = {n50_o, n51_o};
  assign n53_o = t1[14];
  assign n54_o = ~n53_o;
  assign n56_o = {t1, 1'b0};
  assign n57_o = t1s[15:10];
  assign n58_o = t1s[9:0];
  assign n60_o = {1'b0, s0};
  assign n61_o = {n60_o, d1};
  assign n62_o = ~d1;
  assign n63_o = {n61_o, n62_o};
  assign n65_o = {n63_o, 1'b1};
  assign n66_o = t1s_h - u1;
  assign n67_o = d1 ? n66_o : n68_o;
  assign n68_o = t1s_h + u1;
  assign n69_o = t3_h[4:0];
  assign n70_o = {n69_o, t1s_l};
  assign n71_o = {s0, d1};
  assign n72_o = t2[14];
  assign n73_o = ~n72_o;
  assign n75_o = {t2, 1'b0};
  assign n76_o = t2s[15:9];
  assign n77_o = t2s[8:0];
  assign n79_o = {1'b0, s1};
  assign n80_o = {n79_o, d2};
  assign n81_o = ~d2;
  assign n82_o = {n80_o, n81_o};
  assign n84_o = {n82_o, 1'b1};
  assign n85_o = t2s_h - u2;
  assign n86_o = d2 ? n85_o : n87_o;
  assign n87_o = t2s_h + u2;
  assign n88_o = t4_h[5:0];
  assign n89_o = {n88_o, t2s_l};
  assign n90_o = {s1, d2};
  assign n91_o = t3[14];
  assign n92_o = ~n91_o;
  assign n94_o = {t3, 1'b0};
  assign n95_o = t3s[15:8];
  assign n96_o = t3s[7:0];
  assign n98_o = {1'b0, s2};
  assign n99_o = {n98_o, d3};
  assign n100_o = ~d3;
  assign n101_o = {n99_o, n100_o};
  assign n103_o = {n101_o, 1'b1};
  assign n104_o = t3s_h_d1 - u3_d1;
  assign n105_o = d3_d1 ? n104_o : n106_o;
  assign n106_o = t3s_h_d1 + u3_d1;
  assign n107_o = t5_h[6:0];
  assign n108_o = {n107_o, t3s_l_d1};
  assign n109_o = {s2, d3};
  assign n110_o = t4[14];
  assign n111_o = ~n110_o;
  assign n113_o = {t4, 1'b0};
  assign n114_o = t4s[15:7];
  assign n115_o = t4s[6:0];
  assign n117_o = {1'b0, s3_d1};
  assign n118_o = {n117_o, d4};
  assign n119_o = ~d4;
  assign n120_o = {n118_o, n119_o};
  assign n122_o = {n120_o, 1'b1};
  assign n123_o = t4s_h - u4;
  assign n124_o = d4 ? n123_o : n125_o;
  assign n125_o = t4s_h + u4;
  assign n126_o = t6_h[7:0];
  assign n127_o = {n126_o, t4s_l};
  assign n128_o = {s3_d1, d4};
  assign n129_o = t5[14];
  assign n130_o = ~n129_o;
  assign n132_o = {t5, 1'b0};
  assign n133_o = t5s[15:6];
  assign n134_o = t5s[5:0];
  assign n136_o = {1'b0, s4};
  assign n137_o = {n136_o, d5};
  assign n138_o = ~d5;
  assign n139_o = {n137_o, n138_o};
  assign n141_o = {n139_o, 1'b1};
  assign n142_o = t5s_h - u5;
  assign n143_o = d5 ? n142_o : n144_o;
  assign n144_o = t5s_h + u5;
  assign n145_o = t7_h[8:0];
  assign n146_o = {n145_o, t5s_l};
  assign n147_o = {s4, d5};
  assign n148_o = t6[14];
  assign n149_o = ~n148_o;
  assign n151_o = {t6, 1'b0};
  assign n152_o = t6s[15:5];
  assign n153_o = t6s[4:0];
  assign n155_o = {1'b0, s5};
  assign n156_o = {n155_o, d6};
  assign n157_o = ~d6;
  assign n158_o = {n156_o, n157_o};
  assign n160_o = {n158_o, 1'b1};
  assign n161_o = t6s_h - u6;
  assign n162_o = d6 ? n161_o : n163_o;
  assign n163_o = t6s_h + u6;
  assign n164_o = t8_h[9:0];
  assign n165_o = {n164_o, t6s_l};
  assign n166_o = {s5, d6};
  assign n167_o = t7[14];
  assign n168_o = ~n167_o;
  assign n170_o = {t7, 1'b0};
  assign n171_o = t7s[15:4];
  assign n172_o = t7s[3:0];
  assign n174_o = {1'b0, s6};
  assign n175_o = {n174_o, d7};
  assign n176_o = ~d7;
  assign n177_o = {n175_o, n176_o};
  assign n179_o = {n177_o, 1'b1};
  assign n180_o = t7s_h_d1 - u7_d1;
  assign n181_o = d7_d1 ? n180_o : n182_o;
  assign n182_o = t7s_h_d1 + u7_d1;
  assign n183_o = t9_h[10:0];
  assign n184_o = {n183_o, t7s_l_d1};
  assign n185_o = {s6, d7};
  assign n186_o = t8[14];
  assign n187_o = ~n186_o;
  assign n189_o = {t8, 1'b0};
  assign n190_o = t8s[15:3];
  assign n191_o = t8s[2:0];
  assign n193_o = {1'b0, s7_d1};
  assign n194_o = {n193_o, d8};
  assign n195_o = ~d8;
  assign n196_o = {n194_o, n195_o};
  assign n198_o = {n196_o, 1'b1};
  assign n199_o = t8s_h - u8;
  assign n200_o = d8 ? n199_o : n201_o;
  assign n201_o = t8s_h + u8;
  assign n202_o = t10_h[11:0];
  assign n203_o = {n202_o, t8s_l};
  assign n204_o = {s7_d1, d8};
  assign n205_o = t9[14];
  assign n206_o = ~n205_o;
  assign n208_o = {t9, 1'b0};
  assign n209_o = t9s[15:2];
  assign n210_o = t9s[1:0];
  assign n212_o = {1'b0, s8};
  assign n213_o = {n212_o, d9};
  assign n214_o = ~d9;
  assign n215_o = {n213_o, n214_o};
  assign n217_o = {n215_o, 1'b1};
  assign n218_o = t9s_h - u9;
  assign n219_o = d9 ? n218_o : n220_o;
  assign n220_o = t9s_h + u9;
  assign n221_o = t11_h[12:0];
  assign n222_o = {n221_o, t9s_l};
  assign n223_o = {s8, d9};
  assign n224_o = t10[14];
  assign n225_o = ~n224_o;
  assign n227_o = {t10, 1'b0};
  assign n228_o = t10s[15:1];
  assign n229_o = t10s[0];
  assign n231_o = {1'b0, s9};
  assign n232_o = {n231_o, d10};
  assign n233_o = ~d10;
  assign n234_o = {n232_o, n233_o};
  assign n236_o = {n234_o, 1'b1};
  assign n237_o = t10s_h_d1 - u10_d1;
  assign n238_o = d10_d1 ? n237_o : n239_o;
  assign n239_o = t10s_h_d1 + u10_d1;
  assign n240_o = t12_h[13:0];
  assign n241_o = {n240_o, t10s_l_d1};
  assign n242_o = {s9, d10};
  assign n243_o = t11[14];
  assign n244_o = ~n243_o;
  assign n246_o = {t11, 1'b0};
  assign n248_o = {1'b0, s10_d1};
  assign n249_o = {n248_o, d11};
  assign n250_o = ~d11;
  assign n251_o = {n249_o, n250_o};
  assign n253_o = {n251_o, 1'b1};
  assign n254_o = t11s_h - u11;
  assign n255_o = d11 ? n254_o : n256_o;
  assign n256_o = t11s_h + u11;
  assign n257_o = t13_h[14:0];
  assign n258_o = {s10_d1, d11};
  assign n259_o = t12[14];
  assign n260_o = ~n259_o;
  assign n261_o = {s11, d13};
  assign n262_o = mr[11:1];
  assign n263_o = mr[0];
  assign n265_o = {10'b0000000000, round};
  assign n266_o = fr + n265_o;
  assign n267_o = {ern1_d3, frrnd};
  assign n270_o = xsx == 3'b010;
  assign n273_o = xsx == 3'b100;
  assign n276_o = xsx == 3'b000;
  assign n279_o = xsx == 3'b001;
  assign n281_o = {n279_o, n276_o, n273_o, n270_o};
  always @*
    case (n281_o)
      4'b1000: n282_o = 3'b001;
      4'b0100: n282_o = 3'b000;
      4'b0010: n282_o = 3'b100;
      4'b0001: n282_o = 3'b010;
      default: n282_o = 3'b110;
    endcase
  assign n283_o = {xsr_d3, rn2};
  always @(posedge clk)
    n284_q <= ern1;
  always @(posedge clk)
    n285_q <= ern1_d1;
  always @(posedge clk)
    n286_q <= ern1_d2;
  always @(posedge clk)
    n287_q <= d3;
  always @(posedge clk)
    n288_q <= t3s_h;
  always @(posedge clk)
    n289_q <= t3s_l;
  always @(posedge clk)
    n290_q <= u3;
  always @(posedge clk)
    n291_q <= s3;
  always @(posedge clk)
    n292_q <= d7;
  always @(posedge clk)
    n293_q <= t7s_h;
  always @(posedge clk)
    n294_q <= t7s_l;
  always @(posedge clk)
    n295_q <= u7;
  always @(posedge clk)
    n296_q <= s7;
  always @(posedge clk)
    n297_q <= d10;
  always @(posedge clk)
    n298_q <= t10s_h;
  always @(posedge clk)
    n299_q <= t10s_l;
  always @(posedge clk)
    n300_q <= u10;
  always @(posedge clk)
    n301_q <= s10;
  always @(posedge clk)
    n302_q <= xsr;
  always @(posedge clk)
    n303_q <= xsr_d1;
  always @(posedge clk)
    n304_q <= xsr_d2;
endmodule

