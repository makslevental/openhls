module fsqrt#(parameter ID=1)
  (input  clk,
   input  [14:0] X,
   output [14:0] R);
  wire [5:0] fracx;
  wire [5:0] ern0;
  wire [2:0] xsx;
  wire [5:0] ern1;
  wire [5:0] ern1_d1;
  wire [5:0] ern1_d2;
  wire [9:0] fracxnorm;
  wire [1:0] s0;
  wire [9:0] t1;
  wire d1;
  wire [10:0] t1s;
  wire [5:0] t1s_h;
  wire [4:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [9:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [10:0] t2s;
  wire [6:0] t2s_h;
  wire [3:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [9:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [10:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [2:0] t3s_l;
  wire [2:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [9:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [10:0] t4s;
  wire [8:0] t4s_h;
  wire [1:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [9:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [10:0] t5s;
  wire [9:0] t5s_h;
  wire t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [9:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [10:0] t6s;
  wire [10:0] t6s_h;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [9:0] t7;
  wire [7:0] s6;
  wire d8;
  wire [8:0] mr;
  wire [5:0] fr;
  wire [5:0] fr_d1;
  wire round;
  wire round_d1;
  wire [5:0] frrnd;
  wire [11:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [5:0] n16_o;
  wire [4:0] n17_o;
  wire [5:0] n19_o;
  wire [2:0] n20_o;
  wire [5:0] n22_o;
  wire n23_o;
  wire [5:0] n24_o;
  wire [5:0] n25_o;
  wire [6:0] n27_o;
  wire [9:0] n29_o;
  wire n30_o;
  wire n31_o;
  wire [9:0] n32_o;
  wire [7:0] n34_o;
  wire [9:0] n36_o;
  wire [3:0] n38_o;
  wire [3:0] n40_o;
  wire [5:0] n41_o;
  wire [9:0] n42_o;
  wire n43_o;
  wire n44_o;
  wire [10:0] n46_o;
  wire [5:0] n47_o;
  wire [4:0] n48_o;
  wire [2:0] n50_o;
  wire [3:0] n51_o;
  wire n52_o;
  wire [4:0] n53_o;
  wire [5:0] n55_o;
  wire [5:0] n56_o;
  wire [5:0] n57_o;
  wire [5:0] n58_o;
  wire [4:0] n59_o;
  wire [9:0] n60_o;
  wire [2:0] n61_o;
  wire n62_o;
  wire n63_o;
  wire [10:0] n65_o;
  wire [6:0] n66_o;
  wire [3:0] n67_o;
  wire [3:0] n69_o;
  wire [4:0] n70_o;
  wire n71_o;
  wire [5:0] n72_o;
  wire [6:0] n74_o;
  wire [6:0] n75_o;
  wire [6:0] n76_o;
  wire [6:0] n77_o;
  wire [5:0] n78_o;
  wire [9:0] n79_o;
  wire [3:0] n80_o;
  wire n81_o;
  wire n82_o;
  wire [10:0] n84_o;
  wire [7:0] n85_o;
  wire [2:0] n86_o;
  wire [4:0] n88_o;
  wire [5:0] n89_o;
  wire n90_o;
  wire [6:0] n91_o;
  wire [7:0] n93_o;
  wire [7:0] n94_o;
  wire [7:0] n95_o;
  wire [7:0] n96_o;
  wire [6:0] n97_o;
  wire [9:0] n98_o;
  wire [4:0] n99_o;
  wire n100_o;
  wire n101_o;
  wire [10:0] n103_o;
  wire [8:0] n104_o;
  wire [1:0] n105_o;
  wire [5:0] n107_o;
  wire [6:0] n108_o;
  wire n109_o;
  wire [7:0] n110_o;
  wire [8:0] n112_o;
  wire [8:0] n113_o;
  wire [8:0] n114_o;
  wire [8:0] n115_o;
  wire [7:0] n116_o;
  wire [9:0] n117_o;
  wire [5:0] n118_o;
  wire n119_o;
  wire n120_o;
  wire [10:0] n122_o;
  wire [9:0] n123_o;
  wire n124_o;
  wire [6:0] n126_o;
  wire [7:0] n127_o;
  wire n128_o;
  wire [8:0] n129_o;
  wire [9:0] n131_o;
  wire [9:0] n132_o;
  wire [9:0] n133_o;
  wire [9:0] n134_o;
  wire [8:0] n135_o;
  wire [9:0] n136_o;
  wire [6:0] n137_o;
  wire n138_o;
  wire n139_o;
  wire [10:0] n141_o;
  wire [7:0] n143_o;
  wire [8:0] n144_o;
  wire n145_o;
  wire [9:0] n146_o;
  wire [10:0] n148_o;
  wire [10:0] n149_o;
  wire [10:0] n150_o;
  wire [10:0] n151_o;
  wire [9:0] n152_o;
  wire [7:0] n153_o;
  wire n154_o;
  wire n155_o;
  wire [8:0] n156_o;
  wire [5:0] n157_o;
  wire n158_o;
  wire [5:0] n160_o;
  wire [5:0] n161_o;
  wire [11:0] n162_o;
  wire n165_o;
  wire n168_o;
  wire n171_o;
  wire n174_o;
  wire [3:0] n176_o;
  reg [2:0] n177_o;
  wire [14:0] n178_o;
  reg [5:0] n179_q;
  reg [5:0] n180_q;
  reg n181_q;
  reg [7:0] n182_q;
  reg [2:0] n183_q;
  reg [7:0] n184_q;
  reg [4:0] n185_q;
  reg [5:0] n186_q;
  reg n187_q;
  reg [2:0] n188_q;
  reg [2:0] n189_q;
  assign R = n178_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:30:8  */
  assign fracx = n16_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:31:8  */
  assign ern0 = n19_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:32:8  */
  assign xsx = n20_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:33:8  */
  assign ern1 = n25_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:33:14  */
  assign ern1_d1 = n179_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:33:23  */
  assign ern1_d2 = n180_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:34:8  */
  assign fracxnorm = n32_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:36:8  */
  assign t1 = n42_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:37:8  */
  assign d1 = n44_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:38:8  */
  assign t1s = n46_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:39:8  */
  assign t1s_h = n47_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:40:8  */
  assign t1s_l = n48_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:41:8  */
  assign u1 = n55_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:42:8  */
  assign t3_h = n57_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:43:8  */
  assign t2 = n60_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:44:8  */
  assign s1 = n61_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:45:8  */
  assign d2 = n63_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:46:8  */
  assign t2s = n65_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:47:8  */
  assign t2s_h = n66_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:48:8  */
  assign t2s_l = n67_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:49:8  */
  assign u2 = n74_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:50:8  */
  assign t4_h = n76_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:51:8  */
  assign t3 = n79_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:52:8  */
  assign s2 = n80_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:53:8  */
  assign d3 = n82_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:53:12  */
  assign d3_d1 = n181_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:54:8  */
  assign t3s = n84_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:55:8  */
  assign t3s_h = n85_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:55:15  */
  assign t3s_h_d1 = n182_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:56:8  */
  assign t3s_l = n86_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:56:15  */
  assign t3s_l_d1 = n183_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:57:8  */
  assign u3 = n93_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:57:12  */
  assign u3_d1 = n184_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:58:8  */
  assign t5_h = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:59:8  */
  assign t4 = n98_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:60:8  */
  assign s3 = n99_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:60:12  */
  assign s3_d1 = n185_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:61:8  */
  assign d4 = n101_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:62:8  */
  assign t4s = n103_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:63:8  */
  assign t4s_h = n104_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:64:8  */
  assign t4s_l = n105_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:65:8  */
  assign u4 = n112_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:66:8  */
  assign t6_h = n114_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:67:8  */
  assign t5 = n117_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:68:8  */
  assign s4 = n118_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:69:8  */
  assign d5 = n120_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:70:8  */
  assign t5s = n122_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:71:8  */
  assign t5s_h = n123_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:72:8  */
  assign t5s_l = n124_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:73:8  */
  assign u5 = n131_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:74:8  */
  assign t7_h = n133_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:75:8  */
  assign t6 = n136_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:76:8  */
  assign s5 = n137_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:77:8  */
  assign d6 = n139_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:171:16  */
  assign t6s = n141_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:79:8  */
  assign t6s_h = t6s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:80:8  */
  assign u6 = n148_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:81:8  */
  assign t8_h = n150_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:82:8  */
  assign t7 = n152_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:83:8  */
  assign s6 = n153_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:84:8  */
  assign d8 = n155_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:85:8  */
  assign mr = n156_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:86:8  */
  assign fr = n157_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:86:12  */
  assign fr_d1 = n186_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:87:8  */
  assign round = n158_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:87:15  */
  assign round_d1 = n187_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:88:8  */
  assign frrnd = n161_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:89:8  */
  assign rn2 = n162_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:90:8  */
  assign xsr = n177_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:90:13  */
  assign xsr_d1 = n188_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:90:21  */
  assign xsr_d2 = n189_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:108:14  */
  assign n16_o = X[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:109:19  */
  assign n17_o = X[11:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:109:16  */
  assign n19_o = {1'b0, n17_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:110:12  */
  assign n20_o = X[14:12];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:111:17  */
  assign n22_o = ern0 + 6'b001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:111:51  */
  assign n23_o = X[6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:111:48  */
  assign n24_o = {5'b0, n23_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:111:48  */
  assign n25_o = n22_o + n24_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:112:21  */
  assign n27_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:112:29  */
  assign n29_o = {n27_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:112:43  */
  assign n30_o = X[6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:112:47  */
  assign n31_o = ~n30_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:112:37  */
  assign n32_o = n31_o ? n29_o : n36_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:113:15  */
  assign n34_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:113:22  */
  assign n36_o = {n34_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:115:29  */
  assign n38_o = fracxnorm[9:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:115:18  */
  assign n40_o = 4'b0111 + n38_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:115:54  */
  assign n41_o = fracxnorm[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:115:43  */
  assign n42_o = {n40_o, n41_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:119:16  */
  assign n43_o = t1[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:119:10  */
  assign n44_o = ~n43_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:120:14  */
  assign n46_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:121:16  */
  assign n47_o = t1s[10:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:122:16  */
  assign n48_o = t1s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:123:15  */
  assign n50_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:123:20  */
  assign n51_o = {n50_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:123:28  */
  assign n52_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:123:25  */
  assign n53_o = {n51_o, n52_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:123:36  */
  assign n55_o = {n53_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:124:20  */
  assign n56_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:124:25  */
  assign n57_o = d1 ? n56_o : n58_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:125:20  */
  assign n58_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:126:14  */
  assign n59_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:126:27  */
  assign n60_o = {n59_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:127:13  */
  assign n61_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:129:16  */
  assign n62_o = t2[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:129:10  */
  assign n63_o = ~n62_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:130:14  */
  assign n65_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:131:16  */
  assign n66_o = t2s[10:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:132:16  */
  assign n67_o = t2s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:133:15  */
  assign n69_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:133:20  */
  assign n70_o = {n69_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:133:28  */
  assign n71_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:133:25  */
  assign n72_o = {n70_o, n71_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:133:36  */
  assign n74_o = {n72_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:134:20  */
  assign n75_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:134:25  */
  assign n76_o = d2 ? n75_o : n77_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:135:20  */
  assign n77_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:136:14  */
  assign n78_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:136:27  */
  assign n79_o = {n78_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:137:13  */
  assign n80_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:139:16  */
  assign n81_o = t3[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:139:10  */
  assign n82_o = ~n81_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:140:14  */
  assign n84_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:141:16  */
  assign n85_o = t3s[10:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:142:16  */
  assign n86_o = t3s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:143:15  */
  assign n88_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:143:20  */
  assign n89_o = {n88_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:143:28  */
  assign n90_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:143:25  */
  assign n91_o = {n89_o, n90_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:143:36  */
  assign n93_o = {n91_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:144:23  */
  assign n94_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:144:31  */
  assign n95_o = d3_d1 ? n94_o : n96_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:145:23  */
  assign n96_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:146:14  */
  assign n97_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:146:27  */
  assign n98_o = {n97_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:147:13  */
  assign n99_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:149:16  */
  assign n100_o = t4[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:149:10  */
  assign n101_o = ~n100_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:150:14  */
  assign n103_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:151:16  */
  assign n104_o = t4s[10:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:152:16  */
  assign n105_o = t4s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:153:15  */
  assign n107_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:153:23  */
  assign n108_o = {n107_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:153:31  */
  assign n109_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:153:28  */
  assign n110_o = {n108_o, n109_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:153:39  */
  assign n112_o = {n110_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:154:20  */
  assign n113_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:154:25  */
  assign n114_o = d4 ? n113_o : n115_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:155:20  */
  assign n115_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:156:14  */
  assign n116_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:156:27  */
  assign n117_o = {n116_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:157:16  */
  assign n118_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:159:16  */
  assign n119_o = t5[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:159:10  */
  assign n120_o = ~n119_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:160:14  */
  assign n122_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:161:16  */
  assign n123_o = t5s[10:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:162:16  */
  assign n124_o = t5s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:163:15  */
  assign n126_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:163:20  */
  assign n127_o = {n126_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:163:28  */
  assign n128_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:163:25  */
  assign n129_o = {n127_o, n128_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:163:36  */
  assign n131_o = {n129_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:164:20  */
  assign n132_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:164:25  */
  assign n133_o = d5 ? n132_o : n134_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:165:20  */
  assign n134_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:166:14  */
  assign n135_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:166:27  */
  assign n136_o = {n135_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:167:13  */
  assign n137_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:169:16  */
  assign n138_o = t6[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:169:10  */
  assign n139_o = ~n138_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:170:14  */
  assign n141_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:172:15  */
  assign n143_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:172:20  */
  assign n144_o = {n143_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:172:28  */
  assign n145_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:172:25  */
  assign n146_o = {n144_o, n145_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:172:36  */
  assign n148_o = {n146_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:173:20  */
  assign n149_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:173:25  */
  assign n150_o = d6 ? n149_o : n151_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:174:20  */
  assign n151_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:175:14  */
  assign n152_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:176:13  */
  assign n153_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:177:16  */
  assign n154_o = t7[9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:177:10  */
  assign n155_o = ~n154_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:178:13  */
  assign n156_o = {s6, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:179:12  */
  assign n157_o = mr[6:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:180:15  */
  assign n158_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:181:42  */
  assign n160_o = {5'b00000, round_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:181:19  */
  assign n161_o = fr_d1 + n160_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:182:19  */
  assign n162_o = {ern1_d2, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:185:21  */
  assign n165_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:186:21  */
  assign n168_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:187:21  */
  assign n171_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:188:21  */
  assign n174_o = xsx == 3'b001;
  assign n176_o = {n174_o, n171_o, n168_o, n165_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:184:4  */
  always @*
    case (n176_o)
      4'b1000: n177_o = 3'b001;
      4'b0100: n177_o = 3'b000;
      4'b0010: n177_o = 3'b100;
      4'b0001: n177_o = 3'b010;
      default: n177_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:190:16  */
  assign n178_o = {xsr_d2, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n179_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n180_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n181_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n182_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n183_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n184_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n185_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n186_q <= fr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n187_q <= round;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n188_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_6_6.vhdl:94:10  */
  always @(posedge clk)
    n189_q <= xsr_d1;
endmodule

