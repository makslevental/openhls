module selfunction_f300_uid4
    (input wire[8:0] x,
        output wire[2:0] y);
    wire[2:0] y0;
    wire[2:0] y1;
    wire n1127_o;
    wire n1130_o;
    wire n1133_o;
    wire n1136_o;
    wire n1139_o;
    wire n1142_o;
    wire n1145_o;
    wire n1148_o;
    wire n1151_o;
    wire n1154_o;
    wire n1157_o;
    wire n1160_o;
    wire n1163_o;
    wire n1166_o;
    wire n1169_o;
    wire n1172_o;
    wire n1175_o;
    wire n1178_o;
    wire n1181_o;
    wire n1184_o;
    wire n1187_o;
    wire n1190_o;
    wire n1193_o;
    wire n1196_o;
    wire n1199_o;
    wire n1202_o;
    wire n1205_o;
    wire n1208_o;
    wire n1211_o;
    wire n1214_o;
    wire n1217_o;
    wire n1220_o;
    wire n1223_o;
    wire n1226_o;
    wire n1229_o;
    wire n1232_o;
    wire n1235_o;
    wire n1238_o;
    wire n1241_o;
    wire n1244_o;
    wire n1247_o;
    wire n1250_o;
    wire n1253_o;
    wire n1256_o;
    wire n1259_o;
    wire n1262_o;
    wire n1265_o;
    wire n1268_o;
    wire n1271_o;
    wire n1274_o;
    wire n1277_o;
    wire n1280_o;
    wire n1283_o;
    wire n1286_o;
    wire n1289_o;
    wire n1292_o;
    wire n1295_o;
    wire n1298_o;
    wire n1301_o;
    wire n1304_o;
    wire n1307_o;
    wire n1310_o;
    wire n1313_o;
    wire n1316_o;
    wire n1319_o;
    wire n1322_o;
    wire n1325_o;
    wire n1328_o;
    wire n1331_o;
    wire n1334_o;
    wire n1337_o;
    wire n1340_o;
    wire n1343_o;
    wire n1346_o;
    wire n1349_o;
    wire n1352_o;
    wire n1355_o;
    wire n1358_o;
    wire n1361_o;
    wire n1364_o;
    wire n1367_o;
    wire n1370_o;
    wire n1373_o;
    wire n1376_o;
    wire n1379_o;
    wire n1382_o;
    wire n1385_o;
    wire n1388_o;
    wire n1391_o;
    wire n1394_o;
    wire n1397_o;
    wire n1400_o;
    wire n1403_o;
    wire n1406_o;
    wire n1409_o;
    wire n1412_o;
    wire n1415_o;
    wire n1418_o;
    wire n1421_o;
    wire n1424_o;
    wire n1427_o;
    wire n1430_o;
    wire n1433_o;
    wire n1436_o;
    wire n1439_o;
    wire n1442_o;
    wire n1445_o;
    wire n1448_o;
    wire n1451_o;
    wire n1454_o;
    wire n1457_o;
    wire n1460_o;
    wire n1463_o;
    wire n1466_o;
    wire n1469_o;
    wire n1472_o;
    wire n1475_o;
    wire n1478_o;
    wire n1481_o;
    wire n1484_o;
    wire n1487_o;
    wire n1490_o;
    wire n1493_o;
    wire n1496_o;
    wire n1499_o;
    wire n1502_o;
    wire n1505_o;
    wire n1508_o;
    wire n1511_o;
    wire n1514_o;
    wire n1517_o;
    wire n1520_o;
    wire n1523_o;
    wire n1526_o;
    wire n1529_o;
    wire n1532_o;
    wire n1535_o;
    wire n1538_o;
    wire n1541_o;
    wire n1544_o;
    wire n1547_o;
    wire n1550_o;
    wire n1553_o;
    wire n1556_o;
    wire n1559_o;
    wire n1562_o;
    wire n1565_o;
    wire n1568_o;
    wire n1571_o;
    wire n1574_o;
    wire n1577_o;
    wire n1580_o;
    wire n1583_o;
    wire n1586_o;
    wire n1589_o;
    wire n1592_o;
    wire n1595_o;
    wire n1598_o;
    wire n1601_o;
    wire n1604_o;
    wire n1607_o;
    wire n1610_o;
    wire n1613_o;
    wire n1616_o;
    wire n1619_o;
    wire n1622_o;
    wire n1625_o;
    wire n1628_o;
    wire n1631_o;
    wire n1634_o;
    wire n1637_o;
    wire n1640_o;
    wire n1643_o;
    wire n1646_o;
    wire n1649_o;
    wire n1652_o;
    wire n1655_o;
    wire n1658_o;
    wire n1661_o;
    wire n1664_o;
    wire n1667_o;
    wire n1670_o;
    wire n1673_o;
    wire n1676_o;
    wire n1679_o;
    wire n1682_o;
    wire n1685_o;
    wire n1688_o;
    wire n1691_o;
    wire n1694_o;
    wire n1697_o;
    wire n1700_o;
    wire n1703_o;
    wire n1706_o;
    wire n1709_o;
    wire n1712_o;
    wire n1715_o;
    wire n1718_o;
    wire n1721_o;
    wire n1724_o;
    wire n1727_o;
    wire n1730_o;
    wire n1733_o;
    wire n1736_o;
    wire n1739_o;
    wire n1742_o;
    wire n1745_o;
    wire n1748_o;
    wire n1751_o;
    wire n1754_o;
    wire n1757_o;
    wire n1760_o;
    wire n1763_o;
    wire n1766_o;
    wire n1769_o;
    wire n1772_o;
    wire n1775_o;
    wire n1778_o;
    wire n1781_o;
    wire n1784_o;
    wire n1787_o;
    wire n1790_o;
    wire n1793_o;
    wire n1796_o;
    wire n1799_o;
    wire n1802_o;
    wire n1805_o;
    wire n1808_o;
    wire n1811_o;
    wire n1814_o;
    wire n1817_o;
    wire n1820_o;
    wire n1823_o;
    wire n1826_o;
    wire n1829_o;
    wire n1832_o;
    wire n1835_o;
    wire n1838_o;
    wire n1841_o;
    wire n1844_o;
    wire n1847_o;
    wire n1850_o;
    wire n1853_o;
    wire n1856_o;
    wire n1859_o;
    wire n1862_o;
    wire n1865_o;
    wire n1868_o;
    wire n1871_o;
    wire n1874_o;
    wire n1877_o;
    wire n1880_o;
    wire n1883_o;
    wire n1886_o;
    wire n1889_o;
    wire n1892_o;
    wire n1895_o;
    wire n1898_o;
    wire n1901_o;
    wire n1904_o;
    wire n1907_o;
    wire n1910_o;
    wire n1913_o;
    wire n1916_o;
    wire n1919_o;
    wire n1922_o;
    wire n1925_o;
    wire n1928_o;
    wire n1931_o;
    wire n1934_o;
    wire n1937_o;
    wire n1940_o;
    wire n1943_o;
    wire n1946_o;
    wire n1949_o;
    wire n1952_o;
    wire n1955_o;
    wire n1958_o;
    wire n1961_o;
    wire n1964_o;
    wire n1967_o;
    wire n1970_o;
    wire n1973_o;
    wire n1976_o;
    wire n1979_o;
    wire n1982_o;
    wire n1985_o;
    wire n1988_o;
    wire n1991_o;
    wire n1994_o;
    wire n1997_o;
    wire n2000_o;
    wire n2003_o;
    wire n2006_o;
    wire n2009_o;
    wire n2012_o;
    wire n2015_o;
    wire n2018_o;
    wire n2021_o;
    wire n2024_o;
    wire n2027_o;
    wire n2030_o;
    wire n2033_o;
    wire n2036_o;
    wire n2039_o;
    wire n2042_o;
    wire n2045_o;
    wire n2048_o;
    wire n2051_o;
    wire n2054_o;
    wire n2057_o;
    wire n2060_o;
    wire n2063_o;
    wire n2066_o;
    wire n2069_o;
    wire n2072_o;
    wire n2075_o;
    wire n2078_o;
    wire n2081_o;
    wire n2084_o;
    wire n2087_o;
    wire n2090_o;
    wire n2093_o;
    wire n2096_o;
    wire n2099_o;
    wire n2102_o;
    wire n2105_o;
    wire n2108_o;
    wire n2111_o;
    wire n2114_o;
    wire n2117_o;
    wire n2120_o;
    wire n2123_o;
    wire n2126_o;
    wire n2129_o;
    wire n2132_o;
    wire n2135_o;
    wire n2138_o;
    wire n2141_o;
    wire n2144_o;
    wire n2147_o;
    wire n2150_o;
    wire n2153_o;
    wire n2156_o;
    wire n2159_o;
    wire n2162_o;
    wire n2165_o;
    wire n2168_o;
    wire n2171_o;
    wire n2174_o;
    wire n2177_o;
    wire n2180_o;
    wire n2183_o;
    wire n2186_o;
    wire n2189_o;
    wire n2192_o;
    wire n2195_o;
    wire n2198_o;
    wire n2201_o;
    wire n2204_o;
    wire n2207_o;
    wire n2210_o;
    wire n2213_o;
    wire n2216_o;
    wire n2219_o;
    wire n2222_o;
    wire n2225_o;
    wire n2228_o;
    wire n2231_o;
    wire n2234_o;
    wire n2237_o;
    wire n2240_o;
    wire n2243_o;
    wire n2246_o;
    wire n2249_o;
    wire n2252_o;
    wire n2255_o;
    wire n2258_o;
    wire n2261_o;
    wire n2264_o;
    wire n2267_o;
    wire n2270_o;
    wire n2273_o;
    wire n2276_o;
    wire n2279_o;
    wire n2282_o;
    wire n2285_o;
    wire n2288_o;
    wire n2291_o;
    wire n2294_o;
    wire n2297_o;
    wire n2300_o;
    wire n2303_o;
    wire n2306_o;
    wire n2309_o;
    wire n2312_o;
    wire n2315_o;
    wire n2318_o;
    wire n2321_o;
    wire n2324_o;
    wire n2327_o;
    wire n2330_o;
    wire n2333_o;
    wire n2336_o;
    wire n2339_o;
    wire n2342_o;
    wire n2345_o;
    wire n2348_o;
    wire n2351_o;
    wire n2354_o;
    wire n2357_o;
    wire n2360_o;
    wire n2363_o;
    wire n2366_o;
    wire n2369_o;
    wire n2372_o;
    wire n2375_o;
    wire n2378_o;
    wire n2381_o;
    wire n2384_o;
    wire n2387_o;
    wire n2390_o;
    wire n2393_o;
    wire n2396_o;
    wire n2399_o;
    wire n2402_o;
    wire n2405_o;
    wire n2408_o;
    wire n2411_o;
    wire n2414_o;
    wire n2417_o;
    wire n2420_o;
    wire n2423_o;
    wire n2426_o;
    wire n2429_o;
    wire n2432_o;
    wire n2435_o;
    wire n2438_o;
    wire n2441_o;
    wire n2444_o;
    wire n2447_o;
    wire n2450_o;
    wire n2453_o;
    wire n2456_o;
    wire n2459_o;
    wire n2462_o;
    wire n2465_o;
    wire n2468_o;
    wire n2471_o;
    wire n2474_o;
    wire n2477_o;
    wire n2480_o;
    wire n2483_o;
    wire n2486_o;
    wire n2489_o;
    wire n2492_o;
    wire n2495_o;
    wire n2498_o;
    wire n2501_o;
    wire n2504_o;
    wire n2507_o;
    wire n2510_o;
    wire n2513_o;
    wire n2516_o;
    wire n2519_o;
    wire n2522_o;
    wire n2525_o;
    wire n2528_o;
    wire n2531_o;
    wire n2534_o;
    wire n2537_o;
    wire n2540_o;
    wire n2543_o;
    wire n2546_o;
    wire n2549_o;
    wire n2552_o;
    wire n2555_o;
    wire n2558_o;
    wire n2561_o;
    wire n2564_o;
    wire n2567_o;
    wire n2570_o;
    wire n2573_o;
    wire n2576_o;
    wire n2579_o;
    wire n2582_o;
    wire n2585_o;
    wire n2588_o;
    wire n2591_o;
    wire n2594_o;
    wire n2597_o;
    wire n2600_o;
    wire n2603_o;
    wire n2606_o;
    wire n2609_o;
    wire n2612_o;
    wire n2615_o;
    wire n2618_o;
    wire n2621_o;
    wire n2624_o;
    wire n2627_o;
    wire n2630_o;
    wire n2633_o;
    wire n2636_o;
    wire n2639_o;
    wire n2642_o;
    wire n2645_o;
    wire n2648_o;
    wire n2651_o;
    wire n2654_o;
    wire n2657_o;
    wire n2660_o;
    wire[511:0] n2662_o;
    reg[2:0] n2663_o;
    assign y = y1;
    assign y0 = n2663_o; // (signal)
    assign y1 = y0; // (signal)
    assign n1127_o = x == 9'b000000000;
    assign n1130_o = x == 9'b000000001;
    assign n1133_o = x == 9'b000000010;
    assign n1136_o = x == 9'b000000011;
    assign n1139_o = x == 9'b000000100;
    assign n1142_o = x == 9'b000000101;
    assign n1145_o = x == 9'b000000110;
    assign n1148_o = x == 9'b000000111;
    assign n1151_o = x == 9'b000001000;
    assign n1154_o = x == 9'b000001001;
    assign n1157_o = x == 9'b000001010;
    assign n1160_o = x == 9'b000001011;
    assign n1163_o = x == 9'b000001100;
    assign n1166_o = x == 9'b000001101;
    assign n1169_o = x == 9'b000001110;
    assign n1172_o = x == 9'b000001111;
    assign n1175_o = x == 9'b000010000;
    assign n1178_o = x == 9'b000010001;
    assign n1181_o = x == 9'b000010010;
    assign n1184_o = x == 9'b000010011;
    assign n1187_o = x == 9'b000010100;
    assign n1190_o = x == 9'b000010101;
    assign n1193_o = x == 9'b000010110;
    assign n1196_o = x == 9'b000010111;
    assign n1199_o = x == 9'b000011000;
    assign n1202_o = x == 9'b000011001;
    assign n1205_o = x == 9'b000011010;
    assign n1208_o = x == 9'b000011011;
    assign n1211_o = x == 9'b000011100;
    assign n1214_o = x == 9'b000011101;
    assign n1217_o = x == 9'b000011110;
    assign n1220_o = x == 9'b000011111;
    assign n1223_o = x == 9'b000100000;
    assign n1226_o = x == 9'b000100001;
    assign n1229_o = x == 9'b000100010;
    assign n1232_o = x == 9'b000100011;
    assign n1235_o = x == 9'b000100100;
    assign n1238_o = x == 9'b000100101;
    assign n1241_o = x == 9'b000100110;
    assign n1244_o = x == 9'b000100111;
    assign n1247_o = x == 9'b000101000;
    assign n1250_o = x == 9'b000101001;
    assign n1253_o = x == 9'b000101010;
    assign n1256_o = x == 9'b000101011;
    assign n1259_o = x == 9'b000101100;
    assign n1262_o = x == 9'b000101101;
    assign n1265_o = x == 9'b000101110;
    assign n1268_o = x == 9'b000101111;
    assign n1271_o = x == 9'b000110000;
    assign n1274_o = x == 9'b000110001;
    assign n1277_o = x == 9'b000110010;
    assign n1280_o = x == 9'b000110011;
    assign n1283_o = x == 9'b000110100;
    assign n1286_o = x == 9'b000110101;
    assign n1289_o = x == 9'b000110110;
    assign n1292_o = x == 9'b000110111;
    assign n1295_o = x == 9'b000111000;
    assign n1298_o = x == 9'b000111001;
    assign n1301_o = x == 9'b000111010;
    assign n1304_o = x == 9'b000111011;
    assign n1307_o = x == 9'b000111100;
    assign n1310_o = x == 9'b000111101;
    assign n1313_o = x == 9'b000111110;
    assign n1316_o = x == 9'b000111111;
    assign n1319_o = x == 9'b001000000;
    assign n1322_o = x == 9'b001000001;
    assign n1325_o = x == 9'b001000010;
    assign n1328_o = x == 9'b001000011;
    assign n1331_o = x == 9'b001000100;
    assign n1334_o = x == 9'b001000101;
    assign n1337_o = x == 9'b001000110;
    assign n1340_o = x == 9'b001000111;
    assign n1343_o = x == 9'b001001000;
    assign n1346_o = x == 9'b001001001;
    assign n1349_o = x == 9'b001001010;
    assign n1352_o = x == 9'b001001011;
    assign n1355_o = x == 9'b001001100;
    assign n1358_o = x == 9'b001001101;
    assign n1361_o = x == 9'b001001110;
    assign n1364_o = x == 9'b001001111;
    assign n1367_o = x == 9'b001010000;
    assign n1370_o = x == 9'b001010001;
    assign n1373_o = x == 9'b001010010;
    assign n1376_o = x == 9'b001010011;
    assign n1379_o = x == 9'b001010100;
    assign n1382_o = x == 9'b001010101;
    assign n1385_o = x == 9'b001010110;
    assign n1388_o = x == 9'b001010111;
    assign n1391_o = x == 9'b001011000;
    assign n1394_o = x == 9'b001011001;
    assign n1397_o = x == 9'b001011010;
    assign n1400_o = x == 9'b001011011;
    assign n1403_o = x == 9'b001011100;
    assign n1406_o = x == 9'b001011101;
    assign n1409_o = x == 9'b001011110;
    assign n1412_o = x == 9'b001011111;
    assign n1415_o = x == 9'b001100000;
    assign n1418_o = x == 9'b001100001;
    assign n1421_o = x == 9'b001100010;
    assign n1424_o = x == 9'b001100011;
    assign n1427_o = x == 9'b001100100;
    assign n1430_o = x == 9'b001100101;
    assign n1433_o = x == 9'b001100110;
    assign n1436_o = x == 9'b001100111;
    assign n1439_o = x == 9'b001101000;
    assign n1442_o = x == 9'b001101001;
    assign n1445_o = x == 9'b001101010;
    assign n1448_o = x == 9'b001101011;
    assign n1451_o = x == 9'b001101100;
    assign n1454_o = x == 9'b001101101;
    assign n1457_o = x == 9'b001101110;
    assign n1460_o = x == 9'b001101111;
    assign n1463_o = x == 9'b001110000;
    assign n1466_o = x == 9'b001110001;
    assign n1469_o = x == 9'b001110010;
    assign n1472_o = x == 9'b001110011;
    assign n1475_o = x == 9'b001110100;
    assign n1478_o = x == 9'b001110101;
    assign n1481_o = x == 9'b001110110;
    assign n1484_o = x == 9'b001110111;
    assign n1487_o = x == 9'b001111000;
    assign n1490_o = x == 9'b001111001;
    assign n1493_o = x == 9'b001111010;
    assign n1496_o = x == 9'b001111011;
    assign n1499_o = x == 9'b001111100;
    assign n1502_o = x == 9'b001111101;
    assign n1505_o = x == 9'b001111110;
    assign n1508_o = x == 9'b001111111;
    assign n1511_o = x == 9'b010000000;
    assign n1514_o = x == 9'b010000001;
    assign n1517_o = x == 9'b010000010;
    assign n1520_o = x == 9'b010000011;
    assign n1523_o = x == 9'b010000100;
    assign n1526_o = x == 9'b010000101;
    assign n1529_o = x == 9'b010000110;
    assign n1532_o = x == 9'b010000111;
    assign n1535_o = x == 9'b010001000;
    assign n1538_o = x == 9'b010001001;
    assign n1541_o = x == 9'b010001010;
    assign n1544_o = x == 9'b010001011;
    assign n1547_o = x == 9'b010001100;
    assign n1550_o = x == 9'b010001101;
    assign n1553_o = x == 9'b010001110;
    assign n1556_o = x == 9'b010001111;
    assign n1559_o = x == 9'b010010000;
    assign n1562_o = x == 9'b010010001;
    assign n1565_o = x == 9'b010010010;
    assign n1568_o = x == 9'b010010011;
    assign n1571_o = x == 9'b010010100;
    assign n1574_o = x == 9'b010010101;
    assign n1577_o = x == 9'b010010110;
    assign n1580_o = x == 9'b010010111;
    assign n1583_o = x == 9'b010011000;
    assign n1586_o = x == 9'b010011001;
    assign n1589_o = x == 9'b010011010;
    assign n1592_o = x == 9'b010011011;
    assign n1595_o = x == 9'b010011100;
    assign n1598_o = x == 9'b010011101;
    assign n1601_o = x == 9'b010011110;
    assign n1604_o = x == 9'b010011111;
    assign n1607_o = x == 9'b010100000;
    assign n1610_o = x == 9'b010100001;
    assign n1613_o = x == 9'b010100010;
    assign n1616_o = x == 9'b010100011;
    assign n1619_o = x == 9'b010100100;
    assign n1622_o = x == 9'b010100101;
    assign n1625_o = x == 9'b010100110;
    assign n1628_o = x == 9'b010100111;
    assign n1631_o = x == 9'b010101000;
    assign n1634_o = x == 9'b010101001;
    assign n1637_o = x == 9'b010101010;
    assign n1640_o = x == 9'b010101011;
    assign n1643_o = x == 9'b010101100;
    assign n1646_o = x == 9'b010101101;
    assign n1649_o = x == 9'b010101110;
    assign n1652_o = x == 9'b010101111;
    assign n1655_o = x == 9'b010110000;
    assign n1658_o = x == 9'b010110001;
    assign n1661_o = x == 9'b010110010;
    assign n1664_o = x == 9'b010110011;
    assign n1667_o = x == 9'b010110100;
    assign n1670_o = x == 9'b010110101;
    assign n1673_o = x == 9'b010110110;
    assign n1676_o = x == 9'b010110111;
    assign n1679_o = x == 9'b010111000;
    assign n1682_o = x == 9'b010111001;
    assign n1685_o = x == 9'b010111010;
    assign n1688_o = x == 9'b010111011;
    assign n1691_o = x == 9'b010111100;
    assign n1694_o = x == 9'b010111101;
    assign n1697_o = x == 9'b010111110;
    assign n1700_o = x == 9'b010111111;
    assign n1703_o = x == 9'b011000000;
    assign n1706_o = x == 9'b011000001;
    assign n1709_o = x == 9'b011000010;
    assign n1712_o = x == 9'b011000011;
    assign n1715_o = x == 9'b011000100;
    assign n1718_o = x == 9'b011000101;
    assign n1721_o = x == 9'b011000110;
    assign n1724_o = x == 9'b011000111;
    assign n1727_o = x == 9'b011001000;
    assign n1730_o = x == 9'b011001001;
    assign n1733_o = x == 9'b011001010;
    assign n1736_o = x == 9'b011001011;
    assign n1739_o = x == 9'b011001100;
    assign n1742_o = x == 9'b011001101;
    assign n1745_o = x == 9'b011001110;
    assign n1748_o = x == 9'b011001111;
    assign n1751_o = x == 9'b011010000;
    assign n1754_o = x == 9'b011010001;
    assign n1757_o = x == 9'b011010010;
    assign n1760_o = x == 9'b011010011;
    assign n1763_o = x == 9'b011010100;
    assign n1766_o = x == 9'b011010101;
    assign n1769_o = x == 9'b011010110;
    assign n1772_o = x == 9'b011010111;
    assign n1775_o = x == 9'b011011000;
    assign n1778_o = x == 9'b011011001;
    assign n1781_o = x == 9'b011011010;
    assign n1784_o = x == 9'b011011011;
    assign n1787_o = x == 9'b011011100;
    assign n1790_o = x == 9'b011011101;
    assign n1793_o = x == 9'b011011110;
    assign n1796_o = x == 9'b011011111;
    assign n1799_o = x == 9'b011100000;
    assign n1802_o = x == 9'b011100001;
    assign n1805_o = x == 9'b011100010;
    assign n1808_o = x == 9'b011100011;
    assign n1811_o = x == 9'b011100100;
    assign n1814_o = x == 9'b011100101;
    assign n1817_o = x == 9'b011100110;
    assign n1820_o = x == 9'b011100111;
    assign n1823_o = x == 9'b011101000;
    assign n1826_o = x == 9'b011101001;
    assign n1829_o = x == 9'b011101010;
    assign n1832_o = x == 9'b011101011;
    assign n1835_o = x == 9'b011101100;
    assign n1838_o = x == 9'b011101101;
    assign n1841_o = x == 9'b011101110;
    assign n1844_o = x == 9'b011101111;
    assign n1847_o = x == 9'b011110000;
    assign n1850_o = x == 9'b011110001;
    assign n1853_o = x == 9'b011110010;
    assign n1856_o = x == 9'b011110011;
    assign n1859_o = x == 9'b011110100;
    assign n1862_o = x == 9'b011110101;
    assign n1865_o = x == 9'b011110110;
    assign n1868_o = x == 9'b011110111;
    assign n1871_o = x == 9'b011111000;
    assign n1874_o = x == 9'b011111001;
    assign n1877_o = x == 9'b011111010;
    assign n1880_o = x == 9'b011111011;
    assign n1883_o = x == 9'b011111100;
    assign n1886_o = x == 9'b011111101;
    assign n1889_o = x == 9'b011111110;
    assign n1892_o = x == 9'b011111111;
    assign n1895_o = x == 9'b100000000;
    assign n1898_o = x == 9'b100000001;
    assign n1901_o = x == 9'b100000010;
    assign n1904_o = x == 9'b100000011;
    assign n1907_o = x == 9'b100000100;
    assign n1910_o = x == 9'b100000101;
    assign n1913_o = x == 9'b100000110;
    assign n1916_o = x == 9'b100000111;
    assign n1919_o = x == 9'b100001000;
    assign n1922_o = x == 9'b100001001;
    assign n1925_o = x == 9'b100001010;
    assign n1928_o = x == 9'b100001011;
    assign n1931_o = x == 9'b100001100;
    assign n1934_o = x == 9'b100001101;
    assign n1937_o = x == 9'b100001110;
    assign n1940_o = x == 9'b100001111;
    assign n1943_o = x == 9'b100010000;
    assign n1946_o = x == 9'b100010001;
    assign n1949_o = x == 9'b100010010;
    assign n1952_o = x == 9'b100010011;
    assign n1955_o = x == 9'b100010100;
    assign n1958_o = x == 9'b100010101;
    assign n1961_o = x == 9'b100010110;
    assign n1964_o = x == 9'b100010111;
    assign n1967_o = x == 9'b100011000;
    assign n1970_o = x == 9'b100011001;
    assign n1973_o = x == 9'b100011010;
    assign n1976_o = x == 9'b100011011;
    assign n1979_o = x == 9'b100011100;
    assign n1982_o = x == 9'b100011101;
    assign n1985_o = x == 9'b100011110;
    assign n1988_o = x == 9'b100011111;
    assign n1991_o = x == 9'b100100000;
    assign n1994_o = x == 9'b100100001;
    assign n1997_o = x == 9'b100100010;
    assign n2000_o = x == 9'b100100011;
    assign n2003_o = x == 9'b100100100;
    assign n2006_o = x == 9'b100100101;
    assign n2009_o = x == 9'b100100110;
    assign n2012_o = x == 9'b100100111;
    assign n2015_o = x == 9'b100101000;
    assign n2018_o = x == 9'b100101001;
    assign n2021_o = x == 9'b100101010;
    assign n2024_o = x == 9'b100101011;
    assign n2027_o = x == 9'b100101100;
    assign n2030_o = x == 9'b100101101;
    assign n2033_o = x == 9'b100101110;
    assign n2036_o = x == 9'b100101111;
    assign n2039_o = x == 9'b100110000;
    assign n2042_o = x == 9'b100110001;
    assign n2045_o = x == 9'b100110010;
    assign n2048_o = x == 9'b100110011;
    assign n2051_o = x == 9'b100110100;
    assign n2054_o = x == 9'b100110101;
    assign n2057_o = x == 9'b100110110;
    assign n2060_o = x == 9'b100110111;
    assign n2063_o = x == 9'b100111000;
    assign n2066_o = x == 9'b100111001;
    assign n2069_o = x == 9'b100111010;
    assign n2072_o = x == 9'b100111011;
    assign n2075_o = x == 9'b100111100;
    assign n2078_o = x == 9'b100111101;
    assign n2081_o = x == 9'b100111110;
    assign n2084_o = x == 9'b100111111;
    assign n2087_o = x == 9'b101000000;
    assign n2090_o = x == 9'b101000001;
    assign n2093_o = x == 9'b101000010;
    assign n2096_o = x == 9'b101000011;
    assign n2099_o = x == 9'b101000100;
    assign n2102_o = x == 9'b101000101;
    assign n2105_o = x == 9'b101000110;
    assign n2108_o = x == 9'b101000111;
    assign n2111_o = x == 9'b101001000;
    assign n2114_o = x == 9'b101001001;
    assign n2117_o = x == 9'b101001010;
    assign n2120_o = x == 9'b101001011;
    assign n2123_o = x == 9'b101001100;
    assign n2126_o = x == 9'b101001101;
    assign n2129_o = x == 9'b101001110;
    assign n2132_o = x == 9'b101001111;
    assign n2135_o = x == 9'b101010000;
    assign n2138_o = x == 9'b101010001;
    assign n2141_o = x == 9'b101010010;
    assign n2144_o = x == 9'b101010011;
    assign n2147_o = x == 9'b101010100;
    assign n2150_o = x == 9'b101010101;
    assign n2153_o = x == 9'b101010110;
    assign n2156_o = x == 9'b101010111;
    assign n2159_o = x == 9'b101011000;
    assign n2162_o = x == 9'b101011001;
    assign n2165_o = x == 9'b101011010;
    assign n2168_o = x == 9'b101011011;
    assign n2171_o = x == 9'b101011100;
    assign n2174_o = x == 9'b101011101;
    assign n2177_o = x == 9'b101011110;
    assign n2180_o = x == 9'b101011111;
    assign n2183_o = x == 9'b101100000;
    assign n2186_o = x == 9'b101100001;
    assign n2189_o = x == 9'b101100010;
    assign n2192_o = x == 9'b101100011;
    assign n2195_o = x == 9'b101100100;
    assign n2198_o = x == 9'b101100101;
    assign n2201_o = x == 9'b101100110;
    assign n2204_o = x == 9'b101100111;
    assign n2207_o = x == 9'b101101000;
    assign n2210_o = x == 9'b101101001;
    assign n2213_o = x == 9'b101101010;
    assign n2216_o = x == 9'b101101011;
    assign n2219_o = x == 9'b101101100;
    assign n2222_o = x == 9'b101101101;
    assign n2225_o = x == 9'b101101110;
    assign n2228_o = x == 9'b101101111;
    assign n2231_o = x == 9'b101110000;
    assign n2234_o = x == 9'b101110001;
    assign n2237_o = x == 9'b101110010;
    assign n2240_o = x == 9'b101110011;
    assign n2243_o = x == 9'b101110100;
    assign n2246_o = x == 9'b101110101;
    assign n2249_o = x == 9'b101110110;
    assign n2252_o = x == 9'b101110111;
    assign n2255_o = x == 9'b101111000;
    assign n2258_o = x == 9'b101111001;
    assign n2261_o = x == 9'b101111010;
    assign n2264_o = x == 9'b101111011;
    assign n2267_o = x == 9'b101111100;
    assign n2270_o = x == 9'b101111101;
    assign n2273_o = x == 9'b101111110;
    assign n2276_o = x == 9'b101111111;
    assign n2279_o = x == 9'b110000000;
    assign n2282_o = x == 9'b110000001;
    assign n2285_o = x == 9'b110000010;
    assign n2288_o = x == 9'b110000011;
    assign n2291_o = x == 9'b110000100;
    assign n2294_o = x == 9'b110000101;
    assign n2297_o = x == 9'b110000110;
    assign n2300_o = x == 9'b110000111;
    assign n2303_o = x == 9'b110001000;
    assign n2306_o = x == 9'b110001001;
    assign n2309_o = x == 9'b110001010;
    assign n2312_o = x == 9'b110001011;
    assign n2315_o = x == 9'b110001100;
    assign n2318_o = x == 9'b110001101;
    assign n2321_o = x == 9'b110001110;
    assign n2324_o = x == 9'b110001111;
    assign n2327_o = x == 9'b110010000;
    assign n2330_o = x == 9'b110010001;
    assign n2333_o = x == 9'b110010010;
    assign n2336_o = x == 9'b110010011;
    assign n2339_o = x == 9'b110010100;
    assign n2342_o = x == 9'b110010101;
    assign n2345_o = x == 9'b110010110;
    assign n2348_o = x == 9'b110010111;
    assign n2351_o = x == 9'b110011000;
    assign n2354_o = x == 9'b110011001;
    assign n2357_o = x == 9'b110011010;
    assign n2360_o = x == 9'b110011011;
    assign n2363_o = x == 9'b110011100;
    assign n2366_o = x == 9'b110011101;
    assign n2369_o = x == 9'b110011110;
    assign n2372_o = x == 9'b110011111;
    assign n2375_o = x == 9'b110100000;
    assign n2378_o = x == 9'b110100001;
    assign n2381_o = x == 9'b110100010;
    assign n2384_o = x == 9'b110100011;
    assign n2387_o = x == 9'b110100100;
    assign n2390_o = x == 9'b110100101;
    assign n2393_o = x == 9'b110100110;
    assign n2396_o = x == 9'b110100111;
    assign n2399_o = x == 9'b110101000;
    assign n2402_o = x == 9'b110101001;
    assign n2405_o = x == 9'b110101010;
    assign n2408_o = x == 9'b110101011;
    assign n2411_o = x == 9'b110101100;
    assign n2414_o = x == 9'b110101101;
    assign n2417_o = x == 9'b110101110;
    assign n2420_o = x == 9'b110101111;
    assign n2423_o = x == 9'b110110000;
    assign n2426_o = x == 9'b110110001;
    assign n2429_o = x == 9'b110110010;
    assign n2432_o = x == 9'b110110011;
    assign n2435_o = x == 9'b110110100;
    assign n2438_o = x == 9'b110110101;
    assign n2441_o = x == 9'b110110110;
    assign n2444_o = x == 9'b110110111;
    assign n2447_o = x == 9'b110111000;
    assign n2450_o = x == 9'b110111001;
    assign n2453_o = x == 9'b110111010;
    assign n2456_o = x == 9'b110111011;
    assign n2459_o = x == 9'b110111100;
    assign n2462_o = x == 9'b110111101;
    assign n2465_o = x == 9'b110111110;
    assign n2468_o = x == 9'b110111111;
    assign n2471_o = x == 9'b111000000;
    assign n2474_o = x == 9'b111000001;
    assign n2477_o = x == 9'b111000010;
    assign n2480_o = x == 9'b111000011;
    assign n2483_o = x == 9'b111000100;
    assign n2486_o = x == 9'b111000101;
    assign n2489_o = x == 9'b111000110;
    assign n2492_o = x == 9'b111000111;
    assign n2495_o = x == 9'b111001000;
    assign n2498_o = x == 9'b111001001;
    assign n2501_o = x == 9'b111001010;
    assign n2504_o = x == 9'b111001011;
    assign n2507_o = x == 9'b111001100;
    assign n2510_o = x == 9'b111001101;
    assign n2513_o = x == 9'b111001110;
    assign n2516_o = x == 9'b111001111;
    assign n2519_o = x == 9'b111010000;
    assign n2522_o = x == 9'b111010001;
    assign n2525_o = x == 9'b111010010;
    assign n2528_o = x == 9'b111010011;
    assign n2531_o = x == 9'b111010100;
    assign n2534_o = x == 9'b111010101;
    assign n2537_o = x == 9'b111010110;
    assign n2540_o = x == 9'b111010111;
    assign n2543_o = x == 9'b111011000;
    assign n2546_o = x == 9'b111011001;
    assign n2549_o = x == 9'b111011010;
    assign n2552_o = x == 9'b111011011;
    assign n2555_o = x == 9'b111011100;
    assign n2558_o = x == 9'b111011101;
    assign n2561_o = x == 9'b111011110;
    assign n2564_o = x == 9'b111011111;
    assign n2567_o = x == 9'b111100000;
    assign n2570_o = x == 9'b111100001;
    assign n2573_o = x == 9'b111100010;
    assign n2576_o = x == 9'b111100011;
    assign n2579_o = x == 9'b111100100;
    assign n2582_o = x == 9'b111100101;
    assign n2585_o = x == 9'b111100110;
    assign n2588_o = x == 9'b111100111;
    assign n2591_o = x == 9'b111101000;
    assign n2594_o = x == 9'b111101001;
    assign n2597_o = x == 9'b111101010;
    assign n2600_o = x == 9'b111101011;
    assign n2603_o = x == 9'b111101100;
    assign n2606_o = x == 9'b111101101;
    assign n2609_o = x == 9'b111101110;
    assign n2612_o = x == 9'b111101111;
    assign n2615_o = x == 9'b111110000;
    assign n2618_o = x == 9'b111110001;
    assign n2621_o = x == 9'b111110010;
    assign n2624_o = x == 9'b111110011;
    assign n2627_o = x == 9'b111110100;
    assign n2630_o = x == 9'b111110101;
    assign n2633_o = x == 9'b111110110;
    assign n2636_o = x == 9'b111110111;
    assign n2639_o = x == 9'b111111000;
    assign n2642_o = x == 9'b111111001;
    assign n2645_o = x == 9'b111111010;
    assign n2648_o = x == 9'b111111011;
    assign n2651_o = x == 9'b111111100;
    assign n2654_o = x == 9'b111111101;
    assign n2657_o = x == 9'b111111110;
    assign n2660_o = x == 9'b111111111;
    assign n2662_o = {n2660_o, n2657_o, n2654_o, n2651_o, n2648_o, n2645_o, n2642_o, n2639_o, n2636_o, n2633_o, n2630_o, n2627_o, n2624_o, n2621_o, n2618_o, n2615_o, n2612_o, n2609_o, n2606_o, n2603_o, n2600_o, n2597_o, n2594_o, n2591_o, n2588_o, n2585_o, n2582_o, n2579_o, n2576_o, n2573_o, n2570_o, n2567_o, n2564_o, n2561_o, n2558_o, n2555_o, n2552_o, n2549_o, n2546_o, n2543_o, n2540_o, n2537_o, n2534_o, n2531_o, n2528_o, n2525_o, n2522_o, n2519_o, n2516_o, n2513_o, n2510_o, n2507_o, n2504_o, n2501_o, n2498_o, n2495_o, n2492_o, n2489_o, n2486_o, n2483_o, n2480_o, n2477_o, n2474_o, n2471_o, n2468_o, n2465_o, n2462_o, n2459_o, n2456_o, n2453_o, n2450_o, n2447_o, n2444_o, n2441_o, n2438_o, n2435_o, n2432_o, n2429_o, n2426_o, n2423_o, n2420_o, n2417_o, n2414_o, n2411_o, n2408_o, n2405_o, n2402_o, n2399_o, n2396_o, n2393_o, n2390_o, n2387_o, n2384_o, n2381_o, n2378_o, n2375_o, n2372_o, n2369_o, n2366_o, n2363_o, n2360_o, n2357_o, n2354_o, n2351_o, n2348_o, n2345_o, n2342_o, n2339_o, n2336_o, n2333_o, n2330_o, n2327_o, n2324_o, n2321_o, n2318_o, n2315_o, n2312_o, n2309_o, n2306_o, n2303_o, n2300_o, n2297_o, n2294_o, n2291_o, n2288_o, n2285_o, n2282_o, n2279_o, n2276_o, n2273_o, n2270_o, n2267_o, n2264_o, n2261_o, n2258_o, n2255_o, n2252_o, n2249_o, n2246_o, n2243_o, n2240_o, n2237_o, n2234_o, n2231_o, n2228_o, n2225_o, n2222_o, n2219_o, n2216_o, n2213_o, n2210_o, n2207_o, n2204_o, n2201_o, n2198_o, n2195_o, n2192_o, n2189_o, n2186_o, n2183_o, n2180_o, n2177_o, n2174_o, n2171_o, n2168_o, n2165_o, n2162_o, n2159_o, n2156_o, n2153_o, n2150_o, n2147_o, n2144_o, n2141_o, n2138_o, n2135_o, n2132_o, n2129_o, n2126_o, n2123_o, n2120_o, n2117_o, n2114_o, n2111_o, n2108_o, n2105_o, n2102_o, n2099_o, n2096_o, n2093_o, n2090_o, n2087_o, n2084_o, n2081_o, n2078_o, n2075_o, n2072_o, n2069_o, n2066_o, n2063_o, n2060_o, n2057_o, n2054_o, n2051_o, n2048_o, n2045_o, n2042_o, n2039_o, n2036_o, n2033_o, n2030_o, n2027_o, n2024_o, n2021_o, n2018_o, n2015_o, n2012_o, n2009_o, n2006_o, n2003_o, n2000_o, n1997_o, n1994_o, n1991_o, n1988_o, n1985_o, n1982_o, n1979_o, n1976_o, n1973_o, n1970_o, n1967_o, n1964_o, n1961_o, n1958_o, n1955_o, n1952_o, n1949_o, n1946_o, n1943_o, n1940_o, n1937_o, n1934_o, n1931_o, n1928_o, n1925_o, n1922_o, n1919_o, n1916_o, n1913_o, n1910_o, n1907_o, n1904_o, n1901_o, n1898_o, n1895_o, n1892_o, n1889_o, n1886_o, n1883_o, n1880_o, n1877_o, n1874_o, n1871_o, n1868_o, n1865_o, n1862_o, n1859_o, n1856_o, n1853_o, n1850_o, n1847_o, n1844_o, n1841_o, n1838_o, n1835_o, n1832_o, n1829_o, n1826_o, n1823_o, n1820_o, n1817_o, n1814_o, n1811_o, n1808_o, n1805_o, n1802_o, n1799_o, n1796_o, n1793_o, n1790_o, n1787_o, n1784_o, n1781_o, n1778_o, n1775_o, n1772_o, n1769_o, n1766_o, n1763_o, n1760_o, n1757_o, n1754_o, n1751_o, n1748_o, n1745_o, n1742_o, n1739_o, n1736_o, n1733_o, n1730_o, n1727_o, n1724_o, n1721_o, n1718_o, n1715_o, n1712_o, n1709_o, n1706_o, n1703_o, n1700_o, n1697_o, n1694_o, n1691_o, n1688_o, n1685_o, n1682_o, n1679_o, n1676_o, n1673_o, n1670_o, n1667_o, n1664_o, n1661_o, n1658_o, n1655_o, n1652_o, n1649_o, n1646_o, n1643_o, n1640_o, n1637_o, n1634_o, n1631_o, n1628_o, n1625_o, n1622_o, n1619_o, n1616_o, n1613_o, n1610_o, n1607_o, n1604_o, n1601_o, n1598_o, n1595_o, n1592_o, n1589_o, n1586_o, n1583_o, n1580_o, n1577_o, n1574_o, n1571_o, n1568_o, n1565_o, n1562_o, n1559_o, n1556_o, n1553_o, n1550_o, n1547_o, n1544_o, n1541_o, n1538_o, n1535_o, n1532_o, n1529_o, n1526_o, n1523_o, n1520_o, n1517_o, n1514_o, n1511_o, n1508_o, n1505_o, n1502_o, n1499_o, n1496_o, n1493_o, n1490_o, n1487_o, n1484_o, n1481_o, n1478_o, n1475_o, n1472_o, n1469_o, n1466_o, n1463_o, n1460_o, n1457_o, n1454_o, n1451_o, n1448_o, n1445_o, n1442_o, n1439_o, n1436_o, n1433_o, n1430_o, n1427_o, n1424_o, n1421_o, n1418_o, n1415_o, n1412_o, n1409_o, n1406_o, n1403_o, n1400_o, n1397_o, n1394_o, n1391_o, n1388_o, n1385_o, n1382_o, n1379_o, n1376_o, n1373_o, n1370_o, n1367_o, n1364_o, n1361_o, n1358_o, n1355_o, n1352_o, n1349_o, n1346_o, n1343_o, n1340_o, n1337_o, n1334_o, n1331_o, n1328_o, n1325_o, n1322_o, n1319_o, n1316_o, n1313_o, n1310_o, n1307_o, n1304_o, n1301_o, n1298_o, n1295_o, n1292_o, n1289_o, n1286_o, n1283_o, n1280_o, n1277_o, n1274_o, n1271_o, n1268_o, n1265_o, n1262_o, n1259_o, n1256_o, n1253_o, n1250_o, n1247_o, n1244_o, n1241_o, n1238_o, n1235_o, n1232_o, n1229_o, n1226_o, n1223_o, n1220_o, n1217_o, n1214_o, n1211_o, n1208_o, n1205_o, n1202_o, n1199_o, n1196_o, n1193_o, n1190_o, n1187_o, n1184_o, n1181_o, n1178_o, n1175_o, n1172_o, n1169_o, n1166_o, n1163_o, n1160_o, n1157_o, n1154_o, n1151_o, n1148_o, n1145_o, n1142_o, n1139_o, n1136_o, n1133_o, n1130_o, n1127_o};
    always @*
        case (n2662_o)
            512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b111;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b110;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2663_o = 3'b010;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2663_o = 3'b001;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2663_o = 3'b000;
            512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2663_o = 3'b000;
            default: n2663_o = 3'bXXX;
        endcase
endmodule

module fdiv#(parameter ID=1)
    (input wire clk,
        input wire[33:0] X,
        input wire[33:0] Y,
        output wire[33:0] R);
    wire[23:0] fx;
    wire[23:0] fy;
    wire[9:0] expr0;
    wire[9:0] expr0_d1;
    wire[9:0] expr0_d2;
    wire[9:0] expr0_d3;
    wire[9:0] expr0_d4;
    wire[9:0] expr0_d5;
    wire[9:0] expr0_d6;
    wire[9:0] expr0_d7;
    wire[9:0] expr0_d8;
    wire[9:0] expr0_d9;
    wire[9:0] expr0_d10;
    wire[9:0] expr0_d11;
    wire[9:0] expr0_d12;
    wire sr;
    wire sr_d1;
    wire sr_d2;
    wire sr_d3;
    wire sr_d4;
    wire sr_d5;
    wire sr_d6;
    wire sr_d7;
    wire sr_d8;
    wire sr_d9;
    wire sr_d10;
    wire sr_d11;
    wire sr_d12;
    wire[3:0] exnxy;
    wire[1:0] exnr0;
    wire[1:0] exnr0_d1;
    wire[1:0] exnr0_d2;
    wire[1:0] exnr0_d3;
    wire[1:0] exnr0_d4;
    wire[1:0] exnr0_d5;
    wire[1:0] exnr0_d6;
    wire[1:0] exnr0_d7;
    wire[1:0] exnr0_d8;
    wire[1:0] exnr0_d9;
    wire[1:0] exnr0_d10;
    wire[1:0] exnr0_d11;
    wire[1:0] exnr0_d12;
    wire[23:0] d;
    wire[23:0] d_d1;
    wire[23:0] d_d2;
    wire[23:0] d_d3;
    wire[23:0] d_d4;
    wire[23:0] d_d5;
    wire[23:0] d_d6;
    wire[23:0] d_d7;
    wire[23:0] d_d8;
    wire[23:0] d_d9;
    wire[23:0] d_d10;
    wire[23:0] d_d11;
    wire[24:0] psx;
    wire[26:0] betaw14;
    wire[8:0] sel14;
    wire[2:0] q14;
    wire[2:0] q14_copy5;
    wire[26:0] absq14d;
    wire[26:0] w13;
    wire[26:0] betaw13;
    wire[26:0] betaw13_d1;
    wire[8:0] sel13;
    wire[2:0] q13;
    wire[2:0] q13_copy6;
    wire[2:0] q13_copy6_d1;
    wire[26:0] absq13d;
    wire[26:0] w12;
    wire[26:0] betaw12;
    wire[26:0] betaw12_d1;
    wire[8:0] sel12;
    wire[2:0] q12;
    wire[2:0] q12_copy7;
    wire[2:0] q12_copy7_d1;
    wire[26:0] absq12d;
    wire[26:0] w11;
    wire[26:0] betaw11;
    wire[26:0] betaw11_d1;
    wire[8:0] sel11;
    wire[2:0] q11;
    wire[2:0] q11_copy8;
    wire[2:0] q11_copy8_d1;
    wire[26:0] absq11d;
    wire[26:0] w10;
    wire[26:0] betaw10;
    wire[26:0] betaw10_d1;
    wire[8:0] sel10;
    wire[2:0] q10;
    wire[2:0] q10_d1;
    wire[2:0] q10_copy9;
    wire[26:0] absq10d;
    wire[26:0] absq10d_d1;
    wire[26:0] w9;
    wire[26:0] betaw9;
    wire[26:0] betaw9_d1;
    wire[8:0] sel9;
    wire[2:0] q9;
    wire[2:0] q9_d1;
    wire[2:0] q9_copy10;
    wire[26:0] absq9d;
    wire[26:0] absq9d_d1;
    wire[26:0] w8;
    wire[26:0] betaw8;
    wire[26:0] betaw8_d1;
    wire[8:0] sel8;
    wire[2:0] q8;
    wire[2:0] q8_d1;
    wire[2:0] q8_copy11;
    wire[26:0] absq8d;
    wire[26:0] absq8d_d1;
    wire[26:0] w7;
    wire[26:0] betaw7;
    wire[8:0] sel7;
    wire[2:0] q7;
    wire[2:0] q7_copy12;
    wire[26:0] absq7d;
    wire[26:0] w6;
    wire[26:0] betaw6;
    wire[26:0] betaw6_d1;
    wire[8:0] sel6;
    wire[2:0] q6;
    wire[2:0] q6_copy13;
    wire[2:0] q6_copy13_d1;
    wire[26:0] absq6d;
    wire[26:0] w5;
    wire[26:0] betaw5;
    wire[26:0] betaw5_d1;
    wire[8:0] sel5;
    wire[2:0] q5;
    wire[2:0] q5_copy14;
    wire[2:0] q5_copy14_d1;
    wire[26:0] absq5d;
    wire[26:0] w4;
    wire[26:0] betaw4;
    wire[26:0] betaw4_d1;
    wire[8:0] sel4;
    wire[2:0] q4;
    wire[2:0] q4_copy15;
    wire[2:0] q4_copy15_d1;
    wire[26:0] absq4d;
    wire[26:0] w3;
    wire[26:0] betaw3;
    wire[26:0] betaw3_d1;
    wire[8:0] sel3;
    wire[2:0] q3;
    wire[2:0] q3_copy16;
    wire[2:0] q3_copy16_d1;
    wire[26:0] absq3d;
    wire[26:0] w2;
    wire[26:0] betaw2;
    wire[26:0] betaw2_d1;
    wire[8:0] sel2;
    wire[2:0] q2;
    wire[2:0] q2_d1;
    wire[2:0] q2_copy17;
    wire[26:0] absq2d;
    wire[26:0] absq2d_d1;
    wire[26:0] w1;
    wire[26:0] betaw1;
    wire[26:0] betaw1_d1;
    wire[8:0] sel1;
    wire[2:0] q1;
    wire[2:0] q1_d1;
    wire[2:0] q1_copy18;
    wire[26:0] absq1d;
    wire[26:0] absq1d_d1;
    wire[26:0] w0;
    wire[24:0] wfinal;
    wire qm0;
    wire[1:0] qp14;
    wire[1:0] qp14_d1;
    wire[1:0] qp14_d2;
    wire[1:0] qp14_d3;
    wire[1:0] qp14_d4;
    wire[1:0] qp14_d5;
    wire[1:0] qp14_d6;
    wire[1:0] qp14_d7;
    wire[1:0] qp14_d8;
    wire[1:0] qp14_d9;
    wire[1:0] qp14_d10;
    wire[1:0] qp14_d11;
    wire[1:0] qm14;
    wire[1:0] qm14_d1;
    wire[1:0] qm14_d2;
    wire[1:0] qm14_d3;
    wire[1:0] qm14_d4;
    wire[1:0] qm14_d5;
    wire[1:0] qm14_d6;
    wire[1:0] qm14_d7;
    wire[1:0] qm14_d8;
    wire[1:0] qm14_d9;
    wire[1:0] qm14_d10;
    wire[1:0] qm14_d11;
    wire[1:0] qm14_d12;
    wire[1:0] qp13;
    wire[1:0] qp13_d1;
    wire[1:0] qp13_d2;
    wire[1:0] qp13_d3;
    wire[1:0] qp13_d4;
    wire[1:0] qp13_d5;
    wire[1:0] qp13_d6;
    wire[1:0] qp13_d7;
    wire[1:0] qp13_d8;
    wire[1:0] qp13_d9;
    wire[1:0] qp13_d10;
    wire[1:0] qm13;
    wire[1:0] qm13_d1;
    wire[1:0] qm13_d2;
    wire[1:0] qm13_d3;
    wire[1:0] qm13_d4;
    wire[1:0] qm13_d5;
    wire[1:0] qm13_d6;
    wire[1:0] qm13_d7;
    wire[1:0] qm13_d8;
    wire[1:0] qm13_d9;
    wire[1:0] qm13_d10;
    wire[1:0] qm13_d11;
    wire[1:0] qp12;
    wire[1:0] qp12_d1;
    wire[1:0] qp12_d2;
    wire[1:0] qp12_d3;
    wire[1:0] qp12_d4;
    wire[1:0] qp12_d5;
    wire[1:0] qp12_d6;
    wire[1:0] qp12_d7;
    wire[1:0] qp12_d8;
    wire[1:0] qp12_d9;
    wire[1:0] qm12;
    wire[1:0] qm12_d1;
    wire[1:0] qm12_d2;
    wire[1:0] qm12_d3;
    wire[1:0] qm12_d4;
    wire[1:0] qm12_d5;
    wire[1:0] qm12_d6;
    wire[1:0] qm12_d7;
    wire[1:0] qm12_d8;
    wire[1:0] qm12_d9;
    wire[1:0] qm12_d10;
    wire[1:0] qp11;
    wire[1:0] qp11_d1;
    wire[1:0] qp11_d2;
    wire[1:0] qp11_d3;
    wire[1:0] qp11_d4;
    wire[1:0] qp11_d5;
    wire[1:0] qp11_d6;
    wire[1:0] qp11_d7;
    wire[1:0] qp11_d8;
    wire[1:0] qm11;
    wire[1:0] qm11_d1;
    wire[1:0] qm11_d2;
    wire[1:0] qm11_d3;
    wire[1:0] qm11_d4;
    wire[1:0] qm11_d5;
    wire[1:0] qm11_d6;
    wire[1:0] qm11_d7;
    wire[1:0] qm11_d8;
    wire[1:0] qm11_d9;
    wire[1:0] qp10;
    wire[1:0] qp10_d1;
    wire[1:0] qp10_d2;
    wire[1:0] qp10_d3;
    wire[1:0] qp10_d4;
    wire[1:0] qp10_d5;
    wire[1:0] qp10_d6;
    wire[1:0] qp10_d7;
    wire[1:0] qp10_d8;
    wire[1:0] qm10;
    wire[1:0] qm10_d1;
    wire[1:0] qm10_d2;
    wire[1:0] qm10_d3;
    wire[1:0] qm10_d4;
    wire[1:0] qm10_d5;
    wire[1:0] qm10_d6;
    wire[1:0] qm10_d7;
    wire[1:0] qm10_d8;
    wire[1:0] qm10_d9;
    wire[1:0] qp9;
    wire[1:0] qp9_d1;
    wire[1:0] qp9_d2;
    wire[1:0] qp9_d3;
    wire[1:0] qp9_d4;
    wire[1:0] qp9_d5;
    wire[1:0] qp9_d6;
    wire[1:0] qp9_d7;
    wire[1:0] qm9;
    wire[1:0] qm9_d1;
    wire[1:0] qm9_d2;
    wire[1:0] qm9_d3;
    wire[1:0] qm9_d4;
    wire[1:0] qm9_d5;
    wire[1:0] qm9_d6;
    wire[1:0] qm9_d7;
    wire[1:0] qm9_d8;
    wire[1:0] qp8;
    wire[1:0] qp8_d1;
    wire[1:0] qp8_d2;
    wire[1:0] qp8_d3;
    wire[1:0] qp8_d4;
    wire[1:0] qp8_d5;
    wire[1:0] qp8_d6;
    wire[1:0] qm8;
    wire[1:0] qm8_d1;
    wire[1:0] qm8_d2;
    wire[1:0] qm8_d3;
    wire[1:0] qm8_d4;
    wire[1:0] qm8_d5;
    wire[1:0] qm8_d6;
    wire[1:0] qm8_d7;
    wire[1:0] qp7;
    wire[1:0] qp7_d1;
    wire[1:0] qp7_d2;
    wire[1:0] qp7_d3;
    wire[1:0] qp7_d4;
    wire[1:0] qp7_d5;
    wire[1:0] qm7;
    wire[1:0] qm7_d1;
    wire[1:0] qm7_d2;
    wire[1:0] qm7_d3;
    wire[1:0] qm7_d4;
    wire[1:0] qm7_d5;
    wire[1:0] qm7_d6;
    wire[1:0] qp6;
    wire[1:0] qp6_d1;
    wire[1:0] qp6_d2;
    wire[1:0] qp6_d3;
    wire[1:0] qp6_d4;
    wire[1:0] qm6;
    wire[1:0] qm6_d1;
    wire[1:0] qm6_d2;
    wire[1:0] qm6_d3;
    wire[1:0] qm6_d4;
    wire[1:0] qm6_d5;
    wire[1:0] qp5;
    wire[1:0] qp5_d1;
    wire[1:0] qp5_d2;
    wire[1:0] qp5_d3;
    wire[1:0] qm5;
    wire[1:0] qm5_d1;
    wire[1:0] qm5_d2;
    wire[1:0] qm5_d3;
    wire[1:0] qm5_d4;
    wire[1:0] qp4;
    wire[1:0] qp4_d1;
    wire[1:0] qp4_d2;
    wire[1:0] qm4;
    wire[1:0] qm4_d1;
    wire[1:0] qm4_d2;
    wire[1:0] qm4_d3;
    wire[1:0] qp3;
    wire[1:0] qp3_d1;
    wire[1:0] qm3;
    wire[1:0] qm3_d1;
    wire[1:0] qm3_d2;
    wire[1:0] qp2;
    wire[1:0] qp2_d1;
    wire[1:0] qm2;
    wire[1:0] qm2_d1;
    wire[1:0] qm2_d2;
    wire[1:0] qp1;
    wire[1:0] qm1;
    wire[1:0] qm1_d1;
    wire[27:0] qp;
    wire[27:0] qp_d1;
    wire[27:0] qm;
    wire[27:0] quotient;
    wire[25:0] mr;
    wire[23:0] frnorm;
    wire round;
    wire[9:0] expr1;
    wire[32:0] expfrac;
    wire[32:0] expfracr;
    wire[1:0] exnr;
    wire[1:0] exnrfinal;
    wire[22:0] n246_o;
    wire[23:0] n248_o;
    wire[22:0] n249_o;
    wire[23:0] n251_o;
    wire[7:0] n252_o;
    wire[9:0] n254_o;
    wire[7:0] n255_o;
    wire[9:0] n257_o;
    wire[9:0] n258_o;
    wire n259_o;
    wire n260_o;
    wire n261_o;
    wire[1:0] n262_o;
    wire[1:0] n263_o;
    wire[3:0] n264_o;
    wire n267_o;
    wire n270_o;
    wire n272_o;
    wire n273_o;
    wire n275_o;
    wire n276_o;
    wire n279_o;
    wire n281_o;
    wire n282_o;
    wire n284_o;
    wire n285_o;
    wire[2:0] n287_o;
    reg[1:0] n288_o;
    wire[24:0] n290_o;
    wire[26:0] n292_o;
    wire[5:0] n293_o;
    wire[2:0] n294_o;
    wire[8:0] n295_o;
    wire[2:0] selfunctiontable14_n296;
    wire[2:0] selfunctiontable14_y;
    wire[26:0] n300_o;
    wire n302_o;
    wire n304_o;
    wire n305_o;
    wire[25:0] n307_o;
    wire[26:0] n309_o;
    wire n311_o;
    wire n313_o;
    wire n314_o;
    wire[1:0] n316_o;
    reg[26:0] n317_o;
    wire n318_o;
    wire[26:0] n319_o;
    wire n321_o;
    wire[26:0] n322_o;
    reg[26:0] n323_o;
    wire[24:0] n324_o;
    wire[26:0] n326_o;
    wire[5:0] n327_o;
    wire[2:0] n328_o;
    wire[8:0] n329_o;
    wire[2:0] selfunctiontable13_n330;
    wire[2:0] selfunctiontable13_y;
    wire[26:0] n334_o;
    wire n336_o;
    wire n338_o;
    wire n339_o;
    wire[25:0] n341_o;
    wire[26:0] n343_o;
    wire n345_o;
    wire n347_o;
    wire n348_o;
    wire[1:0] n350_o;
    reg[26:0] n351_o;
    wire n352_o;
    wire[26:0] n353_o;
    wire n355_o;
    wire[26:0] n356_o;
    reg[26:0] n357_o;
    wire[24:0] n358_o;
    wire[26:0] n360_o;
    wire[5:0] n361_o;
    wire[2:0] n362_o;
    wire[8:0] n363_o;
    wire[2:0] selfunctiontable12_n364;
    wire[2:0] selfunctiontable12_y;
    wire[26:0] n368_o;
    wire n370_o;
    wire n372_o;
    wire n373_o;
    wire[25:0] n375_o;
    wire[26:0] n377_o;
    wire n379_o;
    wire n381_o;
    wire n382_o;
    wire[1:0] n384_o;
    reg[26:0] n385_o;
    wire n386_o;
    wire[26:0] n387_o;
    wire n389_o;
    wire[26:0] n390_o;
    reg[26:0] n391_o;
    wire[24:0] n392_o;
    wire[26:0] n394_o;
    wire[5:0] n395_o;
    wire[2:0] n396_o;
    wire[8:0] n397_o;
    wire[2:0] selfunctiontable11_n398;
    wire[2:0] selfunctiontable11_y;
    wire[26:0] n402_o;
    wire n404_o;
    wire n406_o;
    wire n407_o;
    wire[25:0] n409_o;
    wire[26:0] n411_o;
    wire n413_o;
    wire n415_o;
    wire n416_o;
    wire[1:0] n418_o;
    reg[26:0] n419_o;
    wire n420_o;
    wire[26:0] n421_o;
    wire n423_o;
    wire[26:0] n424_o;
    reg[26:0] n425_o;
    wire[24:0] n426_o;
    wire[26:0] n428_o;
    wire[5:0] n429_o;
    wire[2:0] n430_o;
    wire[8:0] n431_o;
    wire[2:0] selfunctiontable10_n432;
    wire[2:0] selfunctiontable10_y;
    wire[26:0] n436_o;
    wire n438_o;
    wire n440_o;
    wire n441_o;
    wire[25:0] n443_o;
    wire[26:0] n445_o;
    wire n447_o;
    wire n449_o;
    wire n450_o;
    wire[1:0] n452_o;
    reg[26:0] n453_o;
    wire n454_o;
    wire[26:0] n455_o;
    wire n457_o;
    wire[26:0] n458_o;
    reg[26:0] n459_o;
    wire[24:0] n460_o;
    wire[26:0] n462_o;
    wire[5:0] n463_o;
    wire[2:0] n464_o;
    wire[8:0] n465_o;
    wire[2:0] selfunctiontable9_n466;
    wire[2:0] selfunctiontable9_y;
    wire[26:0] n470_o;
    wire n472_o;
    wire n474_o;
    wire n475_o;
    wire[25:0] n477_o;
    wire[26:0] n479_o;
    wire n481_o;
    wire n483_o;
    wire n484_o;
    wire[1:0] n486_o;
    reg[26:0] n487_o;
    wire n488_o;
    wire[26:0] n489_o;
    wire n491_o;
    wire[26:0] n492_o;
    reg[26:0] n493_o;
    wire[24:0] n494_o;
    wire[26:0] n496_o;
    wire[5:0] n497_o;
    wire[2:0] n498_o;
    wire[8:0] n499_o;
    wire[2:0] selfunctiontable8_n500;
    wire[2:0] selfunctiontable8_y;
    wire[26:0] n504_o;
    wire n506_o;
    wire n508_o;
    wire n509_o;
    wire[25:0] n511_o;
    wire[26:0] n513_o;
    wire n515_o;
    wire n517_o;
    wire n518_o;
    wire[1:0] n520_o;
    reg[26:0] n521_o;
    wire n522_o;
    wire[26:0] n523_o;
    wire n525_o;
    wire[26:0] n526_o;
    reg[26:0] n527_o;
    wire[24:0] n528_o;
    wire[26:0] n530_o;
    wire[5:0] n531_o;
    wire[2:0] n532_o;
    wire[8:0] n533_o;
    wire[2:0] selfunctiontable7_n534;
    wire[2:0] selfunctiontable7_y;
    wire[26:0] n538_o;
    wire n540_o;
    wire n542_o;
    wire n543_o;
    wire[25:0] n545_o;
    wire[26:0] n547_o;
    wire n549_o;
    wire n551_o;
    wire n552_o;
    wire[1:0] n554_o;
    reg[26:0] n555_o;
    wire n556_o;
    wire[26:0] n557_o;
    wire n559_o;
    wire[26:0] n560_o;
    reg[26:0] n561_o;
    wire[24:0] n562_o;
    wire[26:0] n564_o;
    wire[5:0] n565_o;
    wire[2:0] n566_o;
    wire[8:0] n567_o;
    wire[2:0] selfunctiontable6_n568;
    wire[2:0] selfunctiontable6_y;
    wire[26:0] n572_o;
    wire n574_o;
    wire n576_o;
    wire n577_o;
    wire[25:0] n579_o;
    wire[26:0] n581_o;
    wire n583_o;
    wire n585_o;
    wire n586_o;
    wire[1:0] n588_o;
    reg[26:0] n589_o;
    wire n590_o;
    wire[26:0] n591_o;
    wire n593_o;
    wire[26:0] n594_o;
    reg[26:0] n595_o;
    wire[24:0] n596_o;
    wire[26:0] n598_o;
    wire[5:0] n599_o;
    wire[2:0] n600_o;
    wire[8:0] n601_o;
    wire[2:0] selfunctiontable5_n602;
    wire[2:0] selfunctiontable5_y;
    wire[26:0] n606_o;
    wire n608_o;
    wire n610_o;
    wire n611_o;
    wire[25:0] n613_o;
    wire[26:0] n615_o;
    wire n617_o;
    wire n619_o;
    wire n620_o;
    wire[1:0] n622_o;
    reg[26:0] n623_o;
    wire n624_o;
    wire[26:0] n625_o;
    wire n627_o;
    wire[26:0] n628_o;
    reg[26:0] n629_o;
    wire[24:0] n630_o;
    wire[26:0] n632_o;
    wire[5:0] n633_o;
    wire[2:0] n634_o;
    wire[8:0] n635_o;
    wire[2:0] selfunctiontable4_n636;
    wire[2:0] selfunctiontable4_y;
    wire[26:0] n640_o;
    wire n642_o;
    wire n644_o;
    wire n645_o;
    wire[25:0] n647_o;
    wire[26:0] n649_o;
    wire n651_o;
    wire n653_o;
    wire n654_o;
    wire[1:0] n656_o;
    reg[26:0] n657_o;
    wire n658_o;
    wire[26:0] n659_o;
    wire n661_o;
    wire[26:0] n662_o;
    reg[26:0] n663_o;
    wire[24:0] n664_o;
    wire[26:0] n666_o;
    wire[5:0] n667_o;
    wire[2:0] n668_o;
    wire[8:0] n669_o;
    wire[2:0] selfunctiontable3_n670;
    wire[2:0] selfunctiontable3_y;
    wire[26:0] n674_o;
    wire n676_o;
    wire n678_o;
    wire n679_o;
    wire[25:0] n681_o;
    wire[26:0] n683_o;
    wire n685_o;
    wire n687_o;
    wire n688_o;
    wire[1:0] n690_o;
    reg[26:0] n691_o;
    wire n692_o;
    wire[26:0] n693_o;
    wire n695_o;
    wire[26:0] n696_o;
    reg[26:0] n697_o;
    wire[24:0] n698_o;
    wire[26:0] n700_o;
    wire[5:0] n701_o;
    wire[2:0] n702_o;
    wire[8:0] n703_o;
    wire[2:0] selfunctiontable2_n704;
    wire[2:0] selfunctiontable2_y;
    wire[26:0] n708_o;
    wire n710_o;
    wire n712_o;
    wire n713_o;
    wire[25:0] n715_o;
    wire[26:0] n717_o;
    wire n719_o;
    wire n721_o;
    wire n722_o;
    wire[1:0] n724_o;
    reg[26:0] n725_o;
    wire n726_o;
    wire[26:0] n727_o;
    wire n729_o;
    wire[26:0] n730_o;
    reg[26:0] n731_o;
    wire[24:0] n732_o;
    wire[26:0] n734_o;
    wire[5:0] n735_o;
    wire[2:0] n736_o;
    wire[8:0] n737_o;
    wire[2:0] selfunctiontable1_n738;
    wire[2:0] selfunctiontable1_y;
    wire[26:0] n742_o;
    wire n744_o;
    wire n746_o;
    wire n747_o;
    wire[25:0] n749_o;
    wire[26:0] n751_o;
    wire n753_o;
    wire n755_o;
    wire n756_o;
    wire[1:0] n758_o;
    reg[26:0] n759_o;
    wire n760_o;
    wire[26:0] n761_o;
    wire n763_o;
    wire[26:0] n764_o;
    reg[26:0] n765_o;
    wire[24:0] n766_o;
    wire n767_o;
    wire[1:0] n768_o;
    wire n769_o;
    wire[1:0] n771_o;
    wire[1:0] n772_o;
    wire n773_o;
    wire[1:0] n775_o;
    wire[1:0] n776_o;
    wire n777_o;
    wire[1:0] n779_o;
    wire[1:0] n780_o;
    wire n781_o;
    wire[1:0] n783_o;
    wire[1:0] n784_o;
    wire n785_o;
    wire[1:0] n787_o;
    wire[1:0] n788_o;
    wire n789_o;
    wire[1:0] n791_o;
    wire[1:0] n792_o;
    wire n793_o;
    wire[1:0] n795_o;
    wire[1:0] n796_o;
    wire n797_o;
    wire[1:0] n799_o;
    wire[1:0] n800_o;
    wire n801_o;
    wire[1:0] n803_o;
    wire[1:0] n804_o;
    wire n805_o;
    wire[1:0] n807_o;
    wire[1:0] n808_o;
    wire n809_o;
    wire[1:0] n811_o;
    wire[1:0] n812_o;
    wire n813_o;
    wire[1:0] n815_o;
    wire[1:0] n816_o;
    wire n817_o;
    wire[1:0] n819_o;
    wire[1:0] n820_o;
    wire n821_o;
    wire[1:0] n823_o;
    wire[3:0] n824_o;
    wire[5:0] n825_o;
    wire[7:0] n826_o;
    wire[9:0] n827_o;
    wire[11:0] n828_o;
    wire[13:0] n829_o;
    wire[15:0] n830_o;
    wire[17:0] n831_o;
    wire[19:0] n832_o;
    wire[21:0] n833_o;
    wire[23:0] n834_o;
    wire[25:0] n835_o;
    wire[27:0] n836_o;
    wire n837_o;
    wire[2:0] n838_o;
    wire[4:0] n839_o;
    wire[6:0] n840_o;
    wire[8:0] n841_o;
    wire[10:0] n842_o;
    wire[12:0] n843_o;
    wire[14:0] n844_o;
    wire[16:0] n845_o;
    wire[18:0] n846_o;
    wire[20:0] n847_o;
    wire[22:0] n848_o;
    wire[24:0] n849_o;
    wire[26:0] n850_o;
    wire[27:0] n851_o;
    wire[27:0] n852_o;
    wire[25:0] n853_o;
    wire[23:0] n854_o;
    wire n855_o;
    wire[23:0] n856_o;
    wire[23:0] n857_o;
    wire n858_o;
    wire n859_o;
    wire[9:0] n861_o;
    wire[9:0] n862_o;
    wire[22:0] n863_o;
    wire[32:0] n864_o;
    wire[32:0] n866_o;
    wire[32:0] n867_o;
    wire n869_o;
    wire[1:0] n870_o;
    wire[1:0] n872_o;
    wire n874_o;
    wire[1:0] n875_o;
    wire n878_o;
    reg[1:0] n879_o;
    wire[2:0] n880_o;
    wire[30:0] n881_o;
    wire[33:0] n882_o;
    reg[9:0] n883_q;
    reg[9:0] n884_q;
    reg[9:0] n885_q;
    reg[9:0] n886_q;
    reg[9:0] n887_q;
    reg[9:0] n888_q;
    reg[9:0] n889_q;
    reg[9:0] n890_q;
    reg[9:0] n891_q;
    reg[9:0] n892_q;
    reg[9:0] n893_q;
    reg[9:0] n894_q;
    reg n895_q;
    reg n896_q;
    reg n897_q;
    reg n898_q;
    reg n899_q;
    reg n900_q;
    reg n901_q;
    reg n902_q;
    reg n903_q;
    reg n904_q;
    reg n905_q;
    reg n906_q;
    reg[1:0] n907_q;
    reg[1:0] n908_q;
    reg[1:0] n909_q;
    reg[1:0] n910_q;
    reg[1:0] n911_q;
    reg[1:0] n912_q;
    reg[1:0] n913_q;
    reg[1:0] n914_q;
    reg[1:0] n915_q;
    reg[1:0] n916_q;
    reg[1:0] n917_q;
    reg[1:0] n918_q;
    reg[23:0] n919_q;
    reg[23:0] n920_q;
    reg[23:0] n921_q;
    reg[23:0] n922_q;
    reg[23:0] n923_q;
    reg[23:0] n924_q;
    reg[23:0] n925_q;
    reg[23:0] n926_q;
    reg[23:0] n927_q;
    reg[23:0] n928_q;
    reg[23:0] n929_q;
    reg[26:0] n930_q;
    reg[2:0] n931_q;
    reg[26:0] n932_q;
    reg[2:0] n933_q;
    reg[26:0] n934_q;
    reg[2:0] n935_q;
    reg[26:0] n936_q;
    reg[2:0] n937_q;
    reg[26:0] n938_q;
    reg[26:0] n939_q;
    reg[2:0] n940_q;
    reg[26:0] n941_q;
    reg[26:0] n942_q;
    reg[2:0] n943_q;
    reg[26:0] n944_q;
    reg[26:0] n945_q;
    reg[2:0] n946_q;
    reg[26:0] n947_q;
    reg[2:0] n948_q;
    reg[26:0] n949_q;
    reg[2:0] n950_q;
    reg[26:0] n951_q;
    reg[2:0] n952_q;
    reg[26:0] n953_q;
    reg[2:0] n954_q;
    reg[26:0] n955_q;
    reg[26:0] n956_q;
    reg[2:0] n957_q;
    reg[26:0] n958_q;
    reg[1:0] n959_q;
    reg[1:0] n960_q;
    reg[1:0] n961_q;
    reg[1:0] n962_q;
    reg[1:0] n963_q;
    reg[1:0] n964_q;
    reg[1:0] n965_q;
    reg[1:0] n966_q;
    reg[1:0] n967_q;
    reg[1:0] n968_q;
    reg[1:0] n969_q;
    reg[1:0] n970_q;
    reg[1:0] n971_q;
    reg[1:0] n972_q;
    reg[1:0] n973_q;
    reg[1:0] n974_q;
    reg[1:0] n975_q;
    reg[1:0] n976_q;
    reg[1:0] n977_q;
    reg[1:0] n978_q;
    reg[1:0] n979_q;
    reg[1:0] n980_q;
    reg[1:0] n981_q;
    reg[1:0] n982_q;
    reg[1:0] n983_q;
    reg[1:0] n984_q;
    reg[1:0] n985_q;
    reg[1:0] n986_q;
    reg[1:0] n987_q;
    reg[1:0] n988_q;
    reg[1:0] n989_q;
    reg[1:0] n990_q;
    reg[1:0] n991_q;
    reg[1:0] n992_q;
    reg[1:0] n993_q;
    reg[1:0] n994_q;
    reg[1:0] n995_q;
    reg[1:0] n996_q;
    reg[1:0] n997_q;
    reg[1:0] n998_q;
    reg[1:0] n999_q;
    reg[1:0] n1000_q;
    reg[1:0] n1001_q;
    reg[1:0] n1002_q;
    reg[1:0] n1003_q;
    reg[1:0] n1004_q;
    reg[1:0] n1005_q;
    reg[1:0] n1006_q;
    reg[1:0] n1007_q;
    reg[1:0] n1008_q;
    reg[1:0] n1009_q;
    reg[1:0] n1010_q;
    reg[1:0] n1011_q;
    reg[1:0] n1012_q;
    reg[1:0] n1013_q;
    reg[1:0] n1014_q;
    reg[1:0] n1015_q;
    reg[1:0] n1016_q;
    reg[1:0] n1017_q;
    reg[1:0] n1018_q;
    reg[1:0] n1019_q;
    reg[1:0] n1020_q;
    reg[1:0] n1021_q;
    reg[1:0] n1022_q;
    reg[1:0] n1023_q;
    reg[1:0] n1024_q;
    reg[1:0] n1025_q;
    reg[1:0] n1026_q;
    reg[1:0] n1027_q;
    reg[1:0] n1028_q;
    reg[1:0] n1029_q;
    reg[1:0] n1030_q;
    reg[1:0] n1031_q;
    reg[1:0] n1032_q;
    reg[1:0] n1033_q;
    reg[1:0] n1034_q;
    reg[1:0] n1035_q;
    reg[1:0] n1036_q;
    reg[1:0] n1037_q;
    reg[1:0] n1038_q;
    reg[1:0] n1039_q;
    reg[1:0] n1040_q;
    reg[1:0] n1041_q;
    reg[1:0] n1042_q;
    reg[1:0] n1043_q;
    reg[1:0] n1044_q;
    reg[1:0] n1045_q;
    reg[1:0] n1046_q;
    reg[1:0] n1047_q;
    reg[1:0] n1048_q;
    reg[1:0] n1049_q;
    reg[1:0] n1050_q;
    reg[1:0] n1051_q;
    reg[1:0] n1052_q;
    reg[1:0] n1053_q;
    reg[1:0] n1054_q;
    reg[1:0] n1055_q;
    reg[1:0] n1056_q;
    reg[1:0] n1057_q;
    reg[1:0] n1058_q;
    reg[1:0] n1059_q;
    reg[1:0] n1060_q;
    reg[1:0] n1061_q;
    reg[1:0] n1062_q;
    reg[1:0] n1063_q;
    reg[1:0] n1064_q;
    reg[1:0] n1065_q;
    reg[1:0] n1066_q;
    reg[1:0] n1067_q;
    reg[1:0] n1068_q;
    reg[1:0] n1069_q;
    reg[1:0] n1070_q;
    reg[1:0] n1071_q;
    reg[1:0] n1072_q;
    reg[1:0] n1073_q;
    reg[1:0] n1074_q;
    reg[1:0] n1075_q;
    reg[1:0] n1076_q;
    reg[1:0] n1077_q;
    reg[1:0] n1078_q;
    reg[1:0] n1079_q;
    reg[1:0] n1080_q;
    reg[1:0] n1081_q;
    reg[1:0] n1082_q;
    reg[1:0] n1083_q;
    reg[1:0] n1084_q;
    reg[1:0] n1085_q;
    reg[1:0] n1086_q;
    reg[1:0] n1087_q;
    reg[1:0] n1088_q;
    reg[1:0] n1089_q;
    reg[1:0] n1090_q;
    reg[1:0] n1091_q;
    reg[1:0] n1092_q;
    reg[1:0] n1093_q;
    reg[1:0] n1094_q;
    reg[1:0] n1095_q;
    reg[1:0] n1096_q;
    reg[1:0] n1097_q;
    reg[1:0] n1098_q;
    reg[1:0] n1099_q;
    reg[1:0] n1100_q;
    reg[1:0] n1101_q;
    reg[1:0] n1102_q;
    reg[1:0] n1103_q;
    reg[1:0] n1104_q;
    reg[1:0] n1105_q;
    reg[1:0] n1106_q;
    reg[1:0] n1107_q;
    reg[1:0] n1108_q;
    reg[1:0] n1109_q;
    reg[1:0] n1110_q;
    reg[1:0] n1111_q;
    reg[1:0] n1112_q;
    reg[1:0] n1113_q;
    reg[1:0] n1114_q;
    reg[1:0] n1115_q;
    reg[1:0] n1116_q;
    reg[1:0] n1117_q;
    reg[1:0] n1118_q;
    reg[1:0] n1119_q;
    reg[1:0] n1120_q;
    reg[1:0] n1121_q;
    reg[1:0] n1122_q;
    reg[27:0] n1123_q;
    assign R = n882_o;
    assign fx = n248_o; // (signal)
    assign fy = n251_o; // (signal)
    assign expr0 = n258_o; // (signal)
    assign expr0_d1 = n883_q; // (signal)
    assign expr0_d2 = n884_q; // (signal)
    assign expr0_d3 = n885_q; // (signal)
    assign expr0_d4 = n886_q; // (signal)
    assign expr0_d5 = n887_q; // (signal)
    assign expr0_d6 = n888_q; // (signal)
    assign expr0_d7 = n889_q; // (signal)
    assign expr0_d8 = n890_q; // (signal)
    assign expr0_d9 = n891_q; // (signal)
    assign expr0_d10 = n892_q; // (signal)
    assign expr0_d11 = n893_q; // (signal)
    assign expr0_d12 = n894_q; // (signal)
    assign sr = n261_o; // (signal)
    assign sr_d1 = n895_q; // (signal)
    assign sr_d2 = n896_q; // (signal)
    assign sr_d3 = n897_q; // (signal)
    assign sr_d4 = n898_q; // (signal)
    assign sr_d5 = n899_q; // (signal)
    assign sr_d6 = n900_q; // (signal)
    assign sr_d7 = n901_q; // (signal)
    assign sr_d8 = n902_q; // (signal)
    assign sr_d9 = n903_q; // (signal)
    assign sr_d10 = n904_q; // (signal)
    assign sr_d11 = n905_q; // (signal)
    assign sr_d12 = n906_q; // (signal)
    assign exnxy = n264_o; // (signal)
    assign exnr0 = n288_o; // (signal)
    assign exnr0_d1 = n907_q; // (signal)
    assign exnr0_d2 = n908_q; // (signal)
    assign exnr0_d3 = n909_q; // (signal)
    assign exnr0_d4 = n910_q; // (signal)
    assign exnr0_d5 = n911_q; // (signal)
    assign exnr0_d6 = n912_q; // (signal)
    assign exnr0_d7 = n913_q; // (signal)
    assign exnr0_d8 = n914_q; // (signal)
    assign exnr0_d9 = n915_q; // (signal)
    assign exnr0_d10 = n916_q; // (signal)
    assign exnr0_d11 = n917_q; // (signal)
    assign exnr0_d12 = n918_q; // (signal)
    assign d = fy; // (signal)
    assign d_d1 = n919_q; // (signal)
    assign d_d2 = n920_q; // (signal)
    assign d_d3 = n921_q; // (signal)
    assign d_d4 = n922_q; // (signal)
    assign d_d5 = n923_q; // (signal)
    assign d_d6 = n924_q; // (signal)
    assign d_d7 = n925_q; // (signal)
    assign d_d8 = n926_q; // (signal)
    assign d_d9 = n927_q; // (signal)
    assign d_d10 = n928_q; // (signal)
    assign d_d11 = n929_q; // (signal)
    assign psx = n290_o; // (signal)
    assign betaw14 = n292_o; // (signal)
    assign sel14 = n295_o; // (signal)
    assign q14 = q14_copy5; // (signal)
    assign q14_copy5 = selfunctiontable14_n296; // (signal)
    assign absq14d = n317_o; // (signal)
    assign w13 = n323_o; // (signal)
    assign betaw13 = n326_o; // (signal)
    assign betaw13_d1 = n930_q; // (signal)
    assign sel13 = n329_o; // (signal)
    assign q13 = q13_copy6_d1; // (signal)
    assign q13_copy6 = selfunctiontable13_n330; // (signal)
    assign q13_copy6_d1 = n931_q; // (signal)
    assign absq13d = n351_o; // (signal)
    assign w12 = n357_o; // (signal)
    assign betaw12 = n360_o; // (signal)
    assign betaw12_d1 = n932_q; // (signal)
    assign sel12 = n363_o; // (signal)
    assign q12 = q12_copy7_d1; // (signal)
    assign q12_copy7 = selfunctiontable12_n364; // (signal)
    assign q12_copy7_d1 = n933_q; // (signal)
    assign absq12d = n385_o; // (signal)
    assign w11 = n391_o; // (signal)
    assign betaw11 = n394_o; // (signal)
    assign betaw11_d1 = n934_q; // (signal)
    assign sel11 = n397_o; // (signal)
    assign q11 = q11_copy8_d1; // (signal)
    assign q11_copy8 = selfunctiontable11_n398; // (signal)
    assign q11_copy8_d1 = n935_q; // (signal)
    assign absq11d = n419_o; // (signal)
    assign w10 = n425_o; // (signal)
    assign betaw10 = n428_o; // (signal)
    assign betaw10_d1 = n936_q; // (signal)
    assign sel10 = n431_o; // (signal)
    assign q10 = q10_copy9; // (signal)
    assign q10_d1 = n937_q; // (signal)
    assign q10_copy9 = selfunctiontable10_n432; // (signal)
    assign absq10d = n453_o; // (signal)
    assign absq10d_d1 = n938_q; // (signal)
    assign w9 = n459_o; // (signal)
    assign betaw9 = n462_o; // (signal)
    assign betaw9_d1 = n939_q; // (signal)
    assign sel9 = n465_o; // (signal)
    assign q9 = q9_copy10; // (signal)
    assign q9_d1 = n940_q; // (signal)
    assign q9_copy10 = selfunctiontable9_n466; // (signal)
    assign absq9d = n487_o; // (signal)
    assign absq9d_d1 = n941_q; // (signal)
    assign w8 = n493_o; // (signal)
    assign betaw8 = n496_o; // (signal)
    assign betaw8_d1 = n942_q; // (signal)
    assign sel8 = n499_o; // (signal)
    assign q8 = q8_copy11; // (signal)
    assign q8_d1 = n943_q; // (signal)
    assign q8_copy11 = selfunctiontable8_n500; // (signal)
    assign absq8d = n521_o; // (signal)
    assign absq8d_d1 = n944_q; // (signal)
    assign w7 = n527_o; // (signal)
    assign betaw7 = n530_o; // (signal)
    assign sel7 = n533_o; // (signal)
    assign q7 = q7_copy12; // (signal)
    assign q7_copy12 = selfunctiontable7_n534; // (signal)
    assign absq7d = n555_o; // (signal)
    assign w6 = n561_o; // (signal)
    assign betaw6 = n564_o; // (signal)
    assign betaw6_d1 = n945_q; // (signal)
    assign sel6 = n567_o; // (signal)
    assign q6 = q6_copy13_d1; // (signal)
    assign q6_copy13 = selfunctiontable6_n568; // (signal)
    assign q6_copy13_d1 = n946_q; // (signal)
    assign absq6d = n589_o; // (signal)
    assign w5 = n595_o; // (signal)
    assign betaw5 = n598_o; // (signal)
    assign betaw5_d1 = n947_q; // (signal)
    assign sel5 = n601_o; // (signal)
    assign q5 = q5_copy14_d1; // (signal)
    assign q5_copy14 = selfunctiontable5_n602; // (signal)
    assign q5_copy14_d1 = n948_q; // (signal)
    assign absq5d = n623_o; // (signal)
    assign w4 = n629_o; // (signal)
    assign betaw4 = n632_o; // (signal)
    assign betaw4_d1 = n949_q; // (signal)
    assign sel4 = n635_o; // (signal)
    assign q4 = q4_copy15_d1; // (signal)
    assign q4_copy15 = selfunctiontable4_n636; // (signal)
    assign q4_copy15_d1 = n950_q; // (signal)
    assign absq4d = n657_o; // (signal)
    assign w3 = n663_o; // (signal)
    assign betaw3 = n666_o; // (signal)
    assign betaw3_d1 = n951_q; // (signal)
    assign sel3 = n669_o; // (signal)
    assign q3 = q3_copy16_d1; // (signal)
    assign q3_copy16 = selfunctiontable3_n670; // (signal)
    assign q3_copy16_d1 = n952_q; // (signal)
    assign absq3d = n691_o; // (signal)
    assign w2 = n697_o; // (signal)
    assign betaw2 = n700_o; // (signal)
    assign betaw2_d1 = n953_q; // (signal)
    assign sel2 = n703_o; // (signal)
    assign q2 = q2_copy17; // (signal)
    assign q2_d1 = n954_q; // (signal)
    assign q2_copy17 = selfunctiontable2_n704; // (signal)
    assign absq2d = n725_o; // (signal)
    assign absq2d_d1 = n955_q; // (signal)
    assign w1 = n731_o; // (signal)
    assign betaw1 = n734_o; // (signal)
    assign betaw1_d1 = n956_q; // (signal)
    assign sel1 = n737_o; // (signal)
    assign q1 = q1_copy18; // (signal)
    assign q1_d1 = n957_q; // (signal)
    assign q1_copy18 = selfunctiontable1_n738; // (signal)
    assign absq1d = n759_o; // (signal)
    assign absq1d_d1 = n958_q; // (signal)
    assign w0 = n765_o; // (signal)
    assign wfinal = n766_o; // (signal)
    assign qm0 = n767_o; // (signal)
    assign qp14 = n768_o; // (signal)
    assign qp14_d1 = n959_q; // (signal)
    assign qp14_d2 = n960_q; // (signal)
    assign qp14_d3 = n961_q; // (signal)
    assign qp14_d4 = n962_q; // (signal)
    assign qp14_d5 = n963_q; // (signal)
    assign qp14_d6 = n964_q; // (signal)
    assign qp14_d7 = n965_q; // (signal)
    assign qp14_d8 = n966_q; // (signal)
    assign qp14_d9 = n967_q; // (signal)
    assign qp14_d10 = n968_q; // (signal)
    assign qp14_d11 = n969_q; // (signal)
    assign qm14 = n771_o; // (signal)
    assign qm14_d1 = n970_q; // (signal)
    assign qm14_d2 = n971_q; // (signal)
    assign qm14_d3 = n972_q; // (signal)
    assign qm14_d4 = n973_q; // (signal)
    assign qm14_d5 = n974_q; // (signal)
    assign qm14_d6 = n975_q; // (signal)
    assign qm14_d7 = n976_q; // (signal)
    assign qm14_d8 = n977_q; // (signal)
    assign qm14_d9 = n978_q; // (signal)
    assign qm14_d10 = n979_q; // (signal)
    assign qm14_d11 = n980_q; // (signal)
    assign qm14_d12 = n981_q; // (signal)
    assign qp13 = n772_o; // (signal)
    assign qp13_d1 = n982_q; // (signal)
    assign qp13_d2 = n983_q; // (signal)
    assign qp13_d3 = n984_q; // (signal)
    assign qp13_d4 = n985_q; // (signal)
    assign qp13_d5 = n986_q; // (signal)
    assign qp13_d6 = n987_q; // (signal)
    assign qp13_d7 = n988_q; // (signal)
    assign qp13_d8 = n989_q; // (signal)
    assign qp13_d9 = n990_q; // (signal)
    assign qp13_d10 = n991_q; // (signal)
    assign qm13 = n775_o; // (signal)
    assign qm13_d1 = n992_q; // (signal)
    assign qm13_d2 = n993_q; // (signal)
    assign qm13_d3 = n994_q; // (signal)
    assign qm13_d4 = n995_q; // (signal)
    assign qm13_d5 = n996_q; // (signal)
    assign qm13_d6 = n997_q; // (signal)
    assign qm13_d7 = n998_q; // (signal)
    assign qm13_d8 = n999_q; // (signal)
    assign qm13_d9 = n1000_q; // (signal)
    assign qm13_d10 = n1001_q; // (signal)
    assign qm13_d11 = n1002_q; // (signal)
    assign qp12 = n776_o; // (signal)
    assign qp12_d1 = n1003_q; // (signal)
    assign qp12_d2 = n1004_q; // (signal)
    assign qp12_d3 = n1005_q; // (signal)
    assign qp12_d4 = n1006_q; // (signal)
    assign qp12_d5 = n1007_q; // (signal)
    assign qp12_d6 = n1008_q; // (signal)
    assign qp12_d7 = n1009_q; // (signal)
    assign qp12_d8 = n1010_q; // (signal)
    assign qp12_d9 = n1011_q; // (signal)
    assign qm12 = n779_o; // (signal)
    assign qm12_d1 = n1012_q; // (signal)
    assign qm12_d2 = n1013_q; // (signal)
    assign qm12_d3 = n1014_q; // (signal)
    assign qm12_d4 = n1015_q; // (signal)
    assign qm12_d5 = n1016_q; // (signal)
    assign qm12_d6 = n1017_q; // (signal)
    assign qm12_d7 = n1018_q; // (signal)
    assign qm12_d8 = n1019_q; // (signal)
    assign qm12_d9 = n1020_q; // (signal)
    assign qm12_d10 = n1021_q; // (signal)
    assign qp11 = n780_o; // (signal)
    assign qp11_d1 = n1022_q; // (signal)
    assign qp11_d2 = n1023_q; // (signal)
    assign qp11_d3 = n1024_q; // (signal)
    assign qp11_d4 = n1025_q; // (signal)
    assign qp11_d5 = n1026_q; // (signal)
    assign qp11_d6 = n1027_q; // (signal)
    assign qp11_d7 = n1028_q; // (signal)
    assign qp11_d8 = n1029_q; // (signal)
    assign qm11 = n783_o; // (signal)
    assign qm11_d1 = n1030_q; // (signal)
    assign qm11_d2 = n1031_q; // (signal)
    assign qm11_d3 = n1032_q; // (signal)
    assign qm11_d4 = n1033_q; // (signal)
    assign qm11_d5 = n1034_q; // (signal)
    assign qm11_d6 = n1035_q; // (signal)
    assign qm11_d7 = n1036_q; // (signal)
    assign qm11_d8 = n1037_q; // (signal)
    assign qm11_d9 = n1038_q; // (signal)
    assign qp10 = n784_o; // (signal)
    assign qp10_d1 = n1039_q; // (signal)
    assign qp10_d2 = n1040_q; // (signal)
    assign qp10_d3 = n1041_q; // (signal)
    assign qp10_d4 = n1042_q; // (signal)
    assign qp10_d5 = n1043_q; // (signal)
    assign qp10_d6 = n1044_q; // (signal)
    assign qp10_d7 = n1045_q; // (signal)
    assign qp10_d8 = n1046_q; // (signal)
    assign qm10 = n787_o; // (signal)
    assign qm10_d1 = n1047_q; // (signal)
    assign qm10_d2 = n1048_q; // (signal)
    assign qm10_d3 = n1049_q; // (signal)
    assign qm10_d4 = n1050_q; // (signal)
    assign qm10_d5 = n1051_q; // (signal)
    assign qm10_d6 = n1052_q; // (signal)
    assign qm10_d7 = n1053_q; // (signal)
    assign qm10_d8 = n1054_q; // (signal)
    assign qm10_d9 = n1055_q; // (signal)
    assign qp9 = n788_o; // (signal)
    assign qp9_d1 = n1056_q; // (signal)
    assign qp9_d2 = n1057_q; // (signal)
    assign qp9_d3 = n1058_q; // (signal)
    assign qp9_d4 = n1059_q; // (signal)
    assign qp9_d5 = n1060_q; // (signal)
    assign qp9_d6 = n1061_q; // (signal)
    assign qp9_d7 = n1062_q; // (signal)
    assign qm9 = n791_o; // (signal)
    assign qm9_d1 = n1063_q; // (signal)
    assign qm9_d2 = n1064_q; // (signal)
    assign qm9_d3 = n1065_q; // (signal)
    assign qm9_d4 = n1066_q; // (signal)
    assign qm9_d5 = n1067_q; // (signal)
    assign qm9_d6 = n1068_q; // (signal)
    assign qm9_d7 = n1069_q; // (signal)
    assign qm9_d8 = n1070_q; // (signal)
    assign qp8 = n792_o; // (signal)
    assign qp8_d1 = n1071_q; // (signal)
    assign qp8_d2 = n1072_q; // (signal)
    assign qp8_d3 = n1073_q; // (signal)
    assign qp8_d4 = n1074_q; // (signal)
    assign qp8_d5 = n1075_q; // (signal)
    assign qp8_d6 = n1076_q; // (signal)
    assign qm8 = n795_o; // (signal)
    assign qm8_d1 = n1077_q; // (signal)
    assign qm8_d2 = n1078_q; // (signal)
    assign qm8_d3 = n1079_q; // (signal)
    assign qm8_d4 = n1080_q; // (signal)
    assign qm8_d5 = n1081_q; // (signal)
    assign qm8_d6 = n1082_q; // (signal)
    assign qm8_d7 = n1083_q; // (signal)
    assign qp7 = n796_o; // (signal)
    assign qp7_d1 = n1084_q; // (signal)
    assign qp7_d2 = n1085_q; // (signal)
    assign qp7_d3 = n1086_q; // (signal)
    assign qp7_d4 = n1087_q; // (signal)
    assign qp7_d5 = n1088_q; // (signal)
    assign qm7 = n799_o; // (signal)
    assign qm7_d1 = n1089_q; // (signal)
    assign qm7_d2 = n1090_q; // (signal)
    assign qm7_d3 = n1091_q; // (signal)
    assign qm7_d4 = n1092_q; // (signal)
    assign qm7_d5 = n1093_q; // (signal)
    assign qm7_d6 = n1094_q; // (signal)
    assign qp6 = n800_o; // (signal)
    assign qp6_d1 = n1095_q; // (signal)
    assign qp6_d2 = n1096_q; // (signal)
    assign qp6_d3 = n1097_q; // (signal)
    assign qp6_d4 = n1098_q; // (signal)
    assign qm6 = n803_o; // (signal)
    assign qm6_d1 = n1099_q; // (signal)
    assign qm6_d2 = n1100_q; // (signal)
    assign qm6_d3 = n1101_q; // (signal)
    assign qm6_d4 = n1102_q; // (signal)
    assign qm6_d5 = n1103_q; // (signal)
    assign qp5 = n804_o; // (signal)
    assign qp5_d1 = n1104_q; // (signal)
    assign qp5_d2 = n1105_q; // (signal)
    assign qp5_d3 = n1106_q; // (signal)
    assign qm5 = n807_o; // (signal)
    assign qm5_d1 = n1107_q; // (signal)
    assign qm5_d2 = n1108_q; // (signal)
    assign qm5_d3 = n1109_q; // (signal)
    assign qm5_d4 = n1110_q; // (signal)
    assign qp4 = n808_o; // (signal)
    assign qp4_d1 = n1111_q; // (signal)
    assign qp4_d2 = n1112_q; // (signal)
    assign qm4 = n811_o; // (signal)
    assign qm4_d1 = n1113_q; // (signal)
    assign qm4_d2 = n1114_q; // (signal)
    assign qm4_d3 = n1115_q; // (signal)
    assign qp3 = n812_o; // (signal)
    assign qp3_d1 = n1116_q; // (signal)
    assign qm3 = n815_o; // (signal)
    assign qm3_d1 = n1117_q; // (signal)
    assign qm3_d2 = n1118_q; // (signal)
    assign qp2 = n816_o; // (signal)
    assign qp2_d1 = n1119_q; // (signal)
    assign qm2 = n819_o; // (signal)
    assign qm2_d1 = n1120_q; // (signal)
    assign qm2_d2 = n1121_q; // (signal)
    assign qp1 = n820_o; // (signal)
    assign qm1 = n823_o; // (signal)
    assign qm1_d1 = n1122_q; // (signal)
    assign qp = n836_o; // (signal)
    assign qp_d1 = n1123_q; // (signal)
    assign qm = n851_o; // (signal)
    assign quotient = n852_o; // (signal)
    assign mr = n853_o; // (signal)
    assign frnorm = n856_o; // (signal)
    assign round = n858_o; // (signal)
    assign expr1 = n862_o; // (signal)
    assign expfrac = n864_o; // (signal)
    assign expfracr = n867_o; // (signal)
    assign exnr = n870_o; // (signal)
    assign exnrfinal = n879_o; // (signal)
    assign n246_o = X[22:0];
    assign n248_o = {1'b1, n246_o};
    assign n249_o = Y[22:0];
    assign n251_o = {1'b1, n249_o};
    assign n252_o = X[30:23];
    assign n254_o = {2'b00, n252_o};
    assign n255_o = Y[30:23];
    assign n257_o = {2'b00, n255_o};
    assign n258_o = n254_o-n257_o;
    assign n259_o = X[31];
    assign n260_o = Y[31];
    assign n261_o = n259_o ^ n260_o;
    assign n262_o = X[33:32];
    assign n263_o = Y[33:32];
    assign n264_o = {n262_o, n263_o};
    assign n267_o = exnxy == 4'b0101;
    assign n270_o = exnxy == 4'b0001;
    assign n272_o = exnxy == 4'b0010;
    assign n273_o = n270_o | n272_o;
    assign n275_o = exnxy == 4'b0110;
    assign n276_o = n273_o | n275_o;
    assign n279_o = exnxy == 4'b0100;
    assign n281_o = exnxy == 4'b1000;
    assign n282_o = n279_o | n281_o;
    assign n284_o = exnxy == 4'b1001;
    assign n285_o = n282_o | n284_o;
    assign n287_o = {n285_o, n276_o, n267_o};
    always @*
        case (n287_o)
            3'b100: n288_o = 2'b10;
            3'b010: n288_o = 2'b00;
            3'b001: n288_o = 2'b01;
            default: n288_o = 2'b11;
        endcase
    assign n290_o = {1'b0, fx};
    assign n292_o = {2'b00, psx};
    assign n293_o = betaw14[26:21];
    assign n294_o = d[22:20];
    assign n295_o = {n293_o, n294_o};
    assign selfunctiontable14_n296 = selfunctiontable14_y; // (signal)
    selfunction_f300_uid4 selfunctiontable14(
        .x(sel14),
        .y(selfunctiontable14_y));
    assign n300_o = {3'b000, d};
    assign n302_o = q14 == 3'b001;
    assign n304_o = q14 == 3'b111;
    assign n305_o = n302_o | n304_o;
    assign n307_o = {2'b00, d};
    assign n309_o = {n307_o, 1'b0};
    assign n311_o = q14 == 3'b010;
    assign n313_o = q14 == 3'b110;
    assign n314_o = n311_o | n313_o;
    assign n316_o = {n314_o, n305_o};
    always @*
        case (n316_o)
            2'b10: n317_o = n309_o;
            2'b01: n317_o = n300_o;
            default: n317_o = 27'b000000000000000000000000000;
        endcase
    assign n318_o = q14[2];
    assign n319_o = betaw14-absq14d;
    assign n321_o = n318_o == 1'b0;
    assign n322_o = betaw14+absq14d;
    always @*
        case (n321_o)
            1'b1: n323_o = n319_o;
            default: n323_o = n322_o;
        endcase
    assign n324_o = w13[24:0];
    assign n326_o = {n324_o, 2'b00};
    assign n327_o = betaw13[26:21];
    assign n328_o = d[22:20];
    assign n329_o = {n327_o, n328_o};
    assign selfunctiontable13_n330 = selfunctiontable13_y; // (signal)
    selfunction_f300_uid4 selfunctiontable13(
        .x(sel13),
        .y(selfunctiontable13_y));
    assign n334_o = {3'b000, d_d1};
    assign n336_o = q13 == 3'b001;
    assign n338_o = q13 == 3'b111;
    assign n339_o = n336_o | n338_o;
    assign n341_o = {2'b00, d_d1};
    assign n343_o = {n341_o, 1'b0};
    assign n345_o = q13 == 3'b010;
    assign n347_o = q13 == 3'b110;
    assign n348_o = n345_o | n347_o;
    assign n350_o = {n348_o, n339_o};
    always @*
        case (n350_o)
            2'b10: n351_o = n343_o;
            2'b01: n351_o = n334_o;
            default: n351_o = 27'b000000000000000000000000000;
        endcase
    assign n352_o = q13[2];
    assign n353_o = betaw13_d1-absq13d;
    assign n355_o = n352_o == 1'b0;
    assign n356_o = betaw13_d1+absq13d;
    always @*
        case (n355_o)
            1'b1: n357_o = n353_o;
            default: n357_o = n356_o;
        endcase
    assign n358_o = w12[24:0];
    assign n360_o = {n358_o, 2'b00};
    assign n361_o = betaw12[26:21];
    assign n362_o = d_d1[22:20];
    assign n363_o = {n361_o, n362_o};
    assign selfunctiontable12_n364 = selfunctiontable12_y; // (signal)
    selfunction_f300_uid4 selfunctiontable12(
        .x(sel12),
        .y(selfunctiontable12_y));
    assign n368_o = {3'b000, d_d2};
    assign n370_o = q12 == 3'b001;
    assign n372_o = q12 == 3'b111;
    assign n373_o = n370_o | n372_o;
    assign n375_o = {2'b00, d_d2};
    assign n377_o = {n375_o, 1'b0};
    assign n379_o = q12 == 3'b010;
    assign n381_o = q12 == 3'b110;
    assign n382_o = n379_o | n381_o;
    assign n384_o = {n382_o, n373_o};
    always @*
        case (n384_o)
            2'b10: n385_o = n377_o;
            2'b01: n385_o = n368_o;
            default: n385_o = 27'b000000000000000000000000000;
        endcase
    assign n386_o = q12[2];
    assign n387_o = betaw12_d1-absq12d;
    assign n389_o = n386_o == 1'b0;
    assign n390_o = betaw12_d1+absq12d;
    always @*
        case (n389_o)
            1'b1: n391_o = n387_o;
            default: n391_o = n390_o;
        endcase
    assign n392_o = w11[24:0];
    assign n394_o = {n392_o, 2'b00};
    assign n395_o = betaw11[26:21];
    assign n396_o = d_d2[22:20];
    assign n397_o = {n395_o, n396_o};
    assign selfunctiontable11_n398 = selfunctiontable11_y; // (signal)
    selfunction_f300_uid4 selfunctiontable11(
        .x(sel11),
        .y(selfunctiontable11_y));
    assign n402_o = {3'b000, d_d3};
    assign n404_o = q11 == 3'b001;
    assign n406_o = q11 == 3'b111;
    assign n407_o = n404_o | n406_o;
    assign n409_o = {2'b00, d_d3};
    assign n411_o = {n409_o, 1'b0};
    assign n413_o = q11 == 3'b010;
    assign n415_o = q11 == 3'b110;
    assign n416_o = n413_o | n415_o;
    assign n418_o = {n416_o, n407_o};
    always @*
        case (n418_o)
            2'b10: n419_o = n411_o;
            2'b01: n419_o = n402_o;
            default: n419_o = 27'b000000000000000000000000000;
        endcase
    assign n420_o = q11[2];
    assign n421_o = betaw11_d1-absq11d;
    assign n423_o = n420_o == 1'b0;
    assign n424_o = betaw11_d1+absq11d;
    always @*
        case (n423_o)
            1'b1: n425_o = n421_o;
            default: n425_o = n424_o;
        endcase
    assign n426_o = w10[24:0];
    assign n428_o = {n426_o, 2'b00};
    assign n429_o = betaw10[26:21];
    assign n430_o = d_d3[22:20];
    assign n431_o = {n429_o, n430_o};
    assign selfunctiontable10_n432 = selfunctiontable10_y; // (signal)
    selfunction_f300_uid4 selfunctiontable10(
        .x(sel10),
        .y(selfunctiontable10_y));
    assign n436_o = {3'b000, d_d3};
    assign n438_o = q10 == 3'b001;
    assign n440_o = q10 == 3'b111;
    assign n441_o = n438_o | n440_o;
    assign n443_o = {2'b00, d_d3};
    assign n445_o = {n443_o, 1'b0};
    assign n447_o = q10 == 3'b010;
    assign n449_o = q10 == 3'b110;
    assign n450_o = n447_o | n449_o;
    assign n452_o = {n450_o, n441_o};
    always @*
        case (n452_o)
            2'b10: n453_o = n445_o;
            2'b01: n453_o = n436_o;
            default: n453_o = 27'b000000000000000000000000000;
        endcase
    assign n454_o = q10_d1[2];
    assign n455_o = betaw10_d1-absq10d_d1;
    assign n457_o = n454_o == 1'b0;
    assign n458_o = betaw10_d1+absq10d_d1;
    always @*
        case (n457_o)
            1'b1: n459_o = n455_o;
            default: n459_o = n458_o;
        endcase
    assign n460_o = w9[24:0];
    assign n462_o = {n460_o, 2'b00};
    assign n463_o = betaw9[26:21];
    assign n464_o = d_d4[22:20];
    assign n465_o = {n463_o, n464_o};
    assign selfunctiontable9_n466 = selfunctiontable9_y; // (signal)
    selfunction_f300_uid4 selfunctiontable9(
        .x(sel9),
        .y(selfunctiontable9_y));
    assign n470_o = {3'b000, d_d4};
    assign n472_o = q9 == 3'b001;
    assign n474_o = q9 == 3'b111;
    assign n475_o = n472_o | n474_o;
    assign n477_o = {2'b00, d_d4};
    assign n479_o = {n477_o, 1'b0};
    assign n481_o = q9 == 3'b010;
    assign n483_o = q9 == 3'b110;
    assign n484_o = n481_o | n483_o;
    assign n486_o = {n484_o, n475_o};
    always @*
        case (n486_o)
            2'b10: n487_o = n479_o;
            2'b01: n487_o = n470_o;
            default: n487_o = 27'b000000000000000000000000000;
        endcase
    assign n488_o = q9_d1[2];
    assign n489_o = betaw9_d1-absq9d_d1;
    assign n491_o = n488_o == 1'b0;
    assign n492_o = betaw9_d1+absq9d_d1;
    always @*
        case (n491_o)
            1'b1: n493_o = n489_o;
            default: n493_o = n492_o;
        endcase
    assign n494_o = w8[24:0];
    assign n496_o = {n494_o, 2'b00};
    assign n497_o = betaw8[26:21];
    assign n498_o = d_d5[22:20];
    assign n499_o = {n497_o, n498_o};
    assign selfunctiontable8_n500 = selfunctiontable8_y; // (signal)
    selfunction_f300_uid4 selfunctiontable8(
        .x(sel8),
        .y(selfunctiontable8_y));
    assign n504_o = {3'b000, d_d5};
    assign n506_o = q8 == 3'b001;
    assign n508_o = q8 == 3'b111;
    assign n509_o = n506_o | n508_o;
    assign n511_o = {2'b00, d_d5};
    assign n513_o = {n511_o, 1'b0};
    assign n515_o = q8 == 3'b010;
    assign n517_o = q8 == 3'b110;
    assign n518_o = n515_o | n517_o;
    assign n520_o = {n518_o, n509_o};
    always @*
        case (n520_o)
            2'b10: n521_o = n513_o;
            2'b01: n521_o = n504_o;
            default: n521_o = 27'b000000000000000000000000000;
        endcase
    assign n522_o = q8_d1[2];
    assign n523_o = betaw8_d1-absq8d_d1;
    assign n525_o = n522_o == 1'b0;
    assign n526_o = betaw8_d1+absq8d_d1;
    always @*
        case (n525_o)
            1'b1: n527_o = n523_o;
            default: n527_o = n526_o;
        endcase
    assign n528_o = w7[24:0];
    assign n530_o = {n528_o, 2'b00};
    assign n531_o = betaw7[26:21];
    assign n532_o = d_d6[22:20];
    assign n533_o = {n531_o, n532_o};
    assign selfunctiontable7_n534 = selfunctiontable7_y; // (signal)
    selfunction_f300_uid4 selfunctiontable7(
        .x(sel7),
        .y(selfunctiontable7_y));
    assign n538_o = {3'b000, d_d6};
    assign n540_o = q7 == 3'b001;
    assign n542_o = q7 == 3'b111;
    assign n543_o = n540_o | n542_o;
    assign n545_o = {2'b00, d_d6};
    assign n547_o = {n545_o, 1'b0};
    assign n549_o = q7 == 3'b010;
    assign n551_o = q7 == 3'b110;
    assign n552_o = n549_o | n551_o;
    assign n554_o = {n552_o, n543_o};
    always @*
        case (n554_o)
            2'b10: n555_o = n547_o;
            2'b01: n555_o = n538_o;
            default: n555_o = 27'b000000000000000000000000000;
        endcase
    assign n556_o = q7[2];
    assign n557_o = betaw7-absq7d;
    assign n559_o = n556_o == 1'b0;
    assign n560_o = betaw7+absq7d;
    always @*
        case (n559_o)
            1'b1: n561_o = n557_o;
            default: n561_o = n560_o;
        endcase
    assign n562_o = w6[24:0];
    assign n564_o = {n562_o, 2'b00};
    assign n565_o = betaw6[26:21];
    assign n566_o = d_d6[22:20];
    assign n567_o = {n565_o, n566_o};
    assign selfunctiontable6_n568 = selfunctiontable6_y; // (signal)
    selfunction_f300_uid4 selfunctiontable6(
        .x(sel6),
        .y(selfunctiontable6_y));
    assign n572_o = {3'b000, d_d7};
    assign n574_o = q6 == 3'b001;
    assign n576_o = q6 == 3'b111;
    assign n577_o = n574_o | n576_o;
    assign n579_o = {2'b00, d_d7};
    assign n581_o = {n579_o, 1'b0};
    assign n583_o = q6 == 3'b010;
    assign n585_o = q6 == 3'b110;
    assign n586_o = n583_o | n585_o;
    assign n588_o = {n586_o, n577_o};
    always @*
        case (n588_o)
            2'b10: n589_o = n581_o;
            2'b01: n589_o = n572_o;
            default: n589_o = 27'b000000000000000000000000000;
        endcase
    assign n590_o = q6[2];
    assign n591_o = betaw6_d1-absq6d;
    assign n593_o = n590_o == 1'b0;
    assign n594_o = betaw6_d1+absq6d;
    always @*
        case (n593_o)
            1'b1: n595_o = n591_o;
            default: n595_o = n594_o;
        endcase
    assign n596_o = w5[24:0];
    assign n598_o = {n596_o, 2'b00};
    assign n599_o = betaw5[26:21];
    assign n600_o = d_d7[22:20];
    assign n601_o = {n599_o, n600_o};
    assign selfunctiontable5_n602 = selfunctiontable5_y; // (signal)
    selfunction_f300_uid4 selfunctiontable5(
        .x(sel5),
        .y(selfunctiontable5_y));
    assign n606_o = {3'b000, d_d8};
    assign n608_o = q5 == 3'b001;
    assign n610_o = q5 == 3'b111;
    assign n611_o = n608_o | n610_o;
    assign n613_o = {2'b00, d_d8};
    assign n615_o = {n613_o, 1'b0};
    assign n617_o = q5 == 3'b010;
    assign n619_o = q5 == 3'b110;
    assign n620_o = n617_o | n619_o;
    assign n622_o = {n620_o, n611_o};
    always @*
        case (n622_o)
            2'b10: n623_o = n615_o;
            2'b01: n623_o = n606_o;
            default: n623_o = 27'b000000000000000000000000000;
        endcase
    assign n624_o = q5[2];
    assign n625_o = betaw5_d1-absq5d;
    assign n627_o = n624_o == 1'b0;
    assign n628_o = betaw5_d1+absq5d;
    always @*
        case (n627_o)
            1'b1: n629_o = n625_o;
            default: n629_o = n628_o;
        endcase
    assign n630_o = w4[24:0];
    assign n632_o = {n630_o, 2'b00};
    assign n633_o = betaw4[26:21];
    assign n634_o = d_d8[22:20];
    assign n635_o = {n633_o, n634_o};
    assign selfunctiontable4_n636 = selfunctiontable4_y; // (signal)
    selfunction_f300_uid4 selfunctiontable4(
        .x(sel4),
        .y(selfunctiontable4_y));
    assign n640_o = {3'b000, d_d9};
    assign n642_o = q4 == 3'b001;
    assign n644_o = q4 == 3'b111;
    assign n645_o = n642_o | n644_o;
    assign n647_o = {2'b00, d_d9};
    assign n649_o = {n647_o, 1'b0};
    assign n651_o = q4 == 3'b010;
    assign n653_o = q4 == 3'b110;
    assign n654_o = n651_o | n653_o;
    assign n656_o = {n654_o, n645_o};
    always @*
        case (n656_o)
            2'b10: n657_o = n649_o;
            2'b01: n657_o = n640_o;
            default: n657_o = 27'b000000000000000000000000000;
        endcase
    assign n658_o = q4[2];
    assign n659_o = betaw4_d1-absq4d;
    assign n661_o = n658_o == 1'b0;
    assign n662_o = betaw4_d1+absq4d;
    always @*
        case (n661_o)
            1'b1: n663_o = n659_o;
            default: n663_o = n662_o;
        endcase
    assign n664_o = w3[24:0];
    assign n666_o = {n664_o, 2'b00};
    assign n667_o = betaw3[26:21];
    assign n668_o = d_d9[22:20];
    assign n669_o = {n667_o, n668_o};
    assign selfunctiontable3_n670 = selfunctiontable3_y; // (signal)
    selfunction_f300_uid4 selfunctiontable3(
        .x(sel3),
        .y(selfunctiontable3_y));
    assign n674_o = {3'b000, d_d10};
    assign n676_o = q3 == 3'b001;
    assign n678_o = q3 == 3'b111;
    assign n679_o = n676_o | n678_o;
    assign n681_o = {2'b00, d_d10};
    assign n683_o = {n681_o, 1'b0};
    assign n685_o = q3 == 3'b010;
    assign n687_o = q3 == 3'b110;
    assign n688_o = n685_o | n687_o;
    assign n690_o = {n688_o, n679_o};
    always @*
        case (n690_o)
            2'b10: n691_o = n683_o;
            2'b01: n691_o = n674_o;
            default: n691_o = 27'b000000000000000000000000000;
        endcase
    assign n692_o = q3[2];
    assign n693_o = betaw3_d1-absq3d;
    assign n695_o = n692_o == 1'b0;
    assign n696_o = betaw3_d1+absq3d;
    always @*
        case (n695_o)
            1'b1: n697_o = n693_o;
            default: n697_o = n696_o;
        endcase
    assign n698_o = w2[24:0];
    assign n700_o = {n698_o, 2'b00};
    assign n701_o = betaw2[26:21];
    assign n702_o = d_d10[22:20];
    assign n703_o = {n701_o, n702_o};
    assign selfunctiontable2_n704 = selfunctiontable2_y; // (signal)
    selfunction_f300_uid4 selfunctiontable2(
        .x(sel2),
        .y(selfunctiontable2_y));
    assign n708_o = {3'b000, d_d10};
    assign n710_o = q2 == 3'b001;
    assign n712_o = q2 == 3'b111;
    assign n713_o = n710_o | n712_o;
    assign n715_o = {2'b00, d_d10};
    assign n717_o = {n715_o, 1'b0};
    assign n719_o = q2 == 3'b010;
    assign n721_o = q2 == 3'b110;
    assign n722_o = n719_o | n721_o;
    assign n724_o = {n722_o, n713_o};
    always @*
        case (n724_o)
            2'b10: n725_o = n717_o;
            2'b01: n725_o = n708_o;
            default: n725_o = 27'b000000000000000000000000000;
        endcase
    assign n726_o = q2_d1[2];
    assign n727_o = betaw2_d1-absq2d_d1;
    assign n729_o = n726_o == 1'b0;
    assign n730_o = betaw2_d1+absq2d_d1;
    always @*
        case (n729_o)
            1'b1: n731_o = n727_o;
            default: n731_o = n730_o;
        endcase
    assign n732_o = w1[24:0];
    assign n734_o = {n732_o, 2'b00};
    assign n735_o = betaw1[26:21];
    assign n736_o = d_d11[22:20];
    assign n737_o = {n735_o, n736_o};
    assign selfunctiontable1_n738 = selfunctiontable1_y; // (signal)
    selfunction_f300_uid4 selfunctiontable1(
        .x(sel1),
        .y(selfunctiontable1_y));
    assign n742_o = {3'b000, d_d11};
    assign n744_o = q1 == 3'b001;
    assign n746_o = q1 == 3'b111;
    assign n747_o = n744_o | n746_o;
    assign n749_o = {2'b00, d_d11};
    assign n751_o = {n749_o, 1'b0};
    assign n753_o = q1 == 3'b010;
    assign n755_o = q1 == 3'b110;
    assign n756_o = n753_o | n755_o;
    assign n758_o = {n756_o, n747_o};
    always @*
        case (n758_o)
            2'b10: n759_o = n751_o;
            2'b01: n759_o = n742_o;
            default: n759_o = 27'b000000000000000000000000000;
        endcase
    assign n760_o = q1_d1[2];
    assign n761_o = betaw1_d1-absq1d_d1;
    assign n763_o = n760_o == 1'b0;
    assign n764_o = betaw1_d1+absq1d_d1;
    always @*
        case (n763_o)
            1'b1: n765_o = n761_o;
            default: n765_o = n764_o;
        endcase
    assign n766_o = w0[24:0];
    assign n767_o = wfinal[24];
    assign n768_o = q14[1:0];
    assign n769_o = q14[2];
    assign n771_o = {n769_o, 1'b0};
    assign n772_o = q13[1:0];
    assign n773_o = q13[2];
    assign n775_o = {n773_o, 1'b0};
    assign n776_o = q12[1:0];
    assign n777_o = q12[2];
    assign n779_o = {n777_o, 1'b0};
    assign n780_o = q11[1:0];
    assign n781_o = q11[2];
    assign n783_o = {n781_o, 1'b0};
    assign n784_o = q10[1:0];
    assign n785_o = q10[2];
    assign n787_o = {n785_o, 1'b0};
    assign n788_o = q9[1:0];
    assign n789_o = q9[2];
    assign n791_o = {n789_o, 1'b0};
    assign n792_o = q8[1:0];
    assign n793_o = q8[2];
    assign n795_o = {n793_o, 1'b0};
    assign n796_o = q7[1:0];
    assign n797_o = q7[2];
    assign n799_o = {n797_o, 1'b0};
    assign n800_o = q6[1:0];
    assign n801_o = q6[2];
    assign n803_o = {n801_o, 1'b0};
    assign n804_o = q5[1:0];
    assign n805_o = q5[2];
    assign n807_o = {n805_o, 1'b0};
    assign n808_o = q4[1:0];
    assign n809_o = q4[2];
    assign n811_o = {n809_o, 1'b0};
    assign n812_o = q3[1:0];
    assign n813_o = q3[2];
    assign n815_o = {n813_o, 1'b0};
    assign n816_o = q2[1:0];
    assign n817_o = q2[2];
    assign n819_o = {n817_o, 1'b0};
    assign n820_o = q1[1:0];
    assign n821_o = q1[2];
    assign n823_o = {n821_o, 1'b0};
    assign n824_o = {qp14_d11, qp13_d10};
    assign n825_o = {n824_o, qp12_d9};
    assign n826_o = {n825_o, qp11_d8};
    assign n827_o = {n826_o, qp10_d8};
    assign n828_o = {n827_o, qp9_d7};
    assign n829_o = {n828_o, qp8_d6};
    assign n830_o = {n829_o, qp7_d5};
    assign n831_o = {n830_o, qp6_d4};
    assign n832_o = {n831_o, qp5_d3};
    assign n833_o = {n832_o, qp4_d2};
    assign n834_o = {n833_o, qp3_d1};
    assign n835_o = {n834_o, qp2_d1};
    assign n836_o = {n835_o, qp1};
    assign n837_o = qm14_d12[0];
    assign n838_o = {n837_o, qm13_d11};
    assign n839_o = {n838_o, qm12_d10};
    assign n840_o = {n839_o, qm11_d9};
    assign n841_o = {n840_o, qm10_d9};
    assign n842_o = {n841_o, qm9_d8};
    assign n843_o = {n842_o, qm8_d7};
    assign n844_o = {n843_o, qm7_d6};
    assign n845_o = {n844_o, qm6_d5};
    assign n846_o = {n845_o, qm5_d4};
    assign n847_o = {n846_o, qm4_d3};
    assign n848_o = {n847_o, qm3_d2};
    assign n849_o = {n848_o, qm2_d2};
    assign n850_o = {n849_o, qm1_d1};
    assign n851_o = {n850_o, qm0};
    assign n852_o = qp_d1-qm;
    assign n853_o = quotient[26:1];
    assign n854_o = mr[24:1];
    assign n855_o = mr[25];
    assign n856_o = n855_o ? n854_o : n857_o;
    assign n857_o = mr[23:0];
    assign n858_o = frnorm[0];
    assign n859_o = mr[25];
    assign n861_o = {9'b000111111, n859_o};
    assign n862_o = expr0_d12+n861_o;
    assign n863_o = frnorm[23:1];
    assign n864_o = {expr1, n863_o};
    assign n866_o = {32'b00000000000000000000000000000000, round};
    assign n867_o = expfrac+n866_o;
    assign n869_o = expfracr[32];
    assign n870_o = n869_o ? 2'b00 : n875_o;
    assign n872_o = expfracr[32:31];
    assign n874_o = n872_o == 2'b01;
    assign n875_o = n874_o ? 2'b10 : 2'b01;
    assign n878_o = exnr0_d12 == 2'b01;
    always @*
        case (n878_o)
            1'b1: n879_o = exnr;
            default: n879_o = exnr0_d12;
        endcase
    assign n880_o = {exnrfinal, sr_d12};
    assign n881_o = expfracr[30:0];
    assign n882_o = {n880_o, n881_o};
    always @(posedge clk)
        n883_q <= expr0;
    always @(posedge clk)
        n884_q <= expr0_d1;
    always @(posedge clk)
        n885_q <= expr0_d2;
    always @(posedge clk)
        n886_q <= expr0_d3;
    always @(posedge clk)
        n887_q <= expr0_d4;
    always @(posedge clk)
        n888_q <= expr0_d5;
    always @(posedge clk)
        n889_q <= expr0_d6;
    always @(posedge clk)
        n890_q <= expr0_d7;
    always @(posedge clk)
        n891_q <= expr0_d8;
    always @(posedge clk)
        n892_q <= expr0_d9;
    always @(posedge clk)
        n893_q <= expr0_d10;
    always @(posedge clk)
        n894_q <= expr0_d11;
    always @(posedge clk)
        n895_q <= sr;
    always @(posedge clk)
        n896_q <= sr_d1;
    always @(posedge clk)
        n897_q <= sr_d2;
    always @(posedge clk)
        n898_q <= sr_d3;
    always @(posedge clk)
        n899_q <= sr_d4;
    always @(posedge clk)
        n900_q <= sr_d5;
    always @(posedge clk)
        n901_q <= sr_d6;
    always @(posedge clk)
        n902_q <= sr_d7;
    always @(posedge clk)
        n903_q <= sr_d8;
    always @(posedge clk)
        n904_q <= sr_d9;
    always @(posedge clk)
        n905_q <= sr_d10;
    always @(posedge clk)
        n906_q <= sr_d11;
    always @(posedge clk)
        n907_q <= exnr0;
    always @(posedge clk)
        n908_q <= exnr0_d1;
    always @(posedge clk)
        n909_q <= exnr0_d2;
    always @(posedge clk)
        n910_q <= exnr0_d3;
    always @(posedge clk)
        n911_q <= exnr0_d4;
    always @(posedge clk)
        n912_q <= exnr0_d5;
    always @(posedge clk)
        n913_q <= exnr0_d6;
    always @(posedge clk)
        n914_q <= exnr0_d7;
    always @(posedge clk)
        n915_q <= exnr0_d8;
    always @(posedge clk)
        n916_q <= exnr0_d9;
    always @(posedge clk)
        n917_q <= exnr0_d10;
    always @(posedge clk)
        n918_q <= exnr0_d11;
    always @(posedge clk)
        n919_q <= d;
    always @(posedge clk)
        n920_q <= d_d1;
    always @(posedge clk)
        n921_q <= d_d2;
    always @(posedge clk)
        n922_q <= d_d3;
    always @(posedge clk)
        n923_q <= d_d4;
    always @(posedge clk)
        n924_q <= d_d5;
    always @(posedge clk)
        n925_q <= d_d6;
    always @(posedge clk)
        n926_q <= d_d7;
    always @(posedge clk)
        n927_q <= d_d8;
    always @(posedge clk)
        n928_q <= d_d9;
    always @(posedge clk)
        n929_q <= d_d10;
    always @(posedge clk)
        n930_q <= betaw13;
    always @(posedge clk)
        n931_q <= q13_copy6;
    always @(posedge clk)
        n932_q <= betaw12;
    always @(posedge clk)
        n933_q <= q12_copy7;
    always @(posedge clk)
        n934_q <= betaw11;
    always @(posedge clk)
        n935_q <= q11_copy8;
    always @(posedge clk)
        n936_q <= betaw10;
    always @(posedge clk)
        n937_q <= q10;
    always @(posedge clk)
        n938_q <= absq10d;
    always @(posedge clk)
        n939_q <= betaw9;
    always @(posedge clk)
        n940_q <= q9;
    always @(posedge clk)
        n941_q <= absq9d;
    always @(posedge clk)
        n942_q <= betaw8;
    always @(posedge clk)
        n943_q <= q8;
    always @(posedge clk)
        n944_q <= absq8d;
    always @(posedge clk)
        n945_q <= betaw6;
    always @(posedge clk)
        n946_q <= q6_copy13;
    always @(posedge clk)
        n947_q <= betaw5;
    always @(posedge clk)
        n948_q <= q5_copy14;
    always @(posedge clk)
        n949_q <= betaw4;
    always @(posedge clk)
        n950_q <= q4_copy15;
    always @(posedge clk)
        n951_q <= betaw3;
    always @(posedge clk)
        n952_q <= q3_copy16;
    always @(posedge clk)
        n953_q <= betaw2;
    always @(posedge clk)
        n954_q <= q2;
    always @(posedge clk)
        n955_q <= absq2d;
    always @(posedge clk)
        n956_q <= betaw1;
    always @(posedge clk)
        n957_q <= q1;
    always @(posedge clk)
        n958_q <= absq1d;
    always @(posedge clk)
        n959_q <= qp14;
    always @(posedge clk)
        n960_q <= qp14_d1;
    always @(posedge clk)
        n961_q <= qp14_d2;
    always @(posedge clk)
        n962_q <= qp14_d3;
    always @(posedge clk)
        n963_q <= qp14_d4;
    always @(posedge clk)
        n964_q <= qp14_d5;
    always @(posedge clk)
        n965_q <= qp14_d6;
    always @(posedge clk)
        n966_q <= qp14_d7;
    always @(posedge clk)
        n967_q <= qp14_d8;
    always @(posedge clk)
        n968_q <= qp14_d9;
    always @(posedge clk)
        n969_q <= qp14_d10;
    always @(posedge clk)
        n970_q <= qm14;
    always @(posedge clk)
        n971_q <= qm14_d1;
    always @(posedge clk)
        n972_q <= qm14_d2;
    always @(posedge clk)
        n973_q <= qm14_d3;
    always @(posedge clk)
        n974_q <= qm14_d4;
    always @(posedge clk)
        n975_q <= qm14_d5;
    always @(posedge clk)
        n976_q <= qm14_d6;
    always @(posedge clk)
        n977_q <= qm14_d7;
    always @(posedge clk)
        n978_q <= qm14_d8;
    always @(posedge clk)
        n979_q <= qm14_d9;
    always @(posedge clk)
        n980_q <= qm14_d10;
    always @(posedge clk)
        n981_q <= qm14_d11;
    always @(posedge clk)
        n982_q <= qp13;
    always @(posedge clk)
        n983_q <= qp13_d1;
    always @(posedge clk)
        n984_q <= qp13_d2;
    always @(posedge clk)
        n985_q <= qp13_d3;
    always @(posedge clk)
        n986_q <= qp13_d4;
    always @(posedge clk)
        n987_q <= qp13_d5;
    always @(posedge clk)
        n988_q <= qp13_d6;
    always @(posedge clk)
        n989_q <= qp13_d7;
    always @(posedge clk)
        n990_q <= qp13_d8;
    always @(posedge clk)
        n991_q <= qp13_d9;
    always @(posedge clk)
        n992_q <= qm13;
    always @(posedge clk)
        n993_q <= qm13_d1;
    always @(posedge clk)
        n994_q <= qm13_d2;
    always @(posedge clk)
        n995_q <= qm13_d3;
    always @(posedge clk)
        n996_q <= qm13_d4;
    always @(posedge clk)
        n997_q <= qm13_d5;
    always @(posedge clk)
        n998_q <= qm13_d6;
    always @(posedge clk)
        n999_q <= qm13_d7;
    always @(posedge clk)
        n1000_q <= qm13_d8;
    always @(posedge clk)
        n1001_q <= qm13_d9;
    always @(posedge clk)
        n1002_q <= qm13_d10;
    always @(posedge clk)
        n1003_q <= qp12;
    always @(posedge clk)
        n1004_q <= qp12_d1;
    always @(posedge clk)
        n1005_q <= qp12_d2;
    always @(posedge clk)
        n1006_q <= qp12_d3;
    always @(posedge clk)
        n1007_q <= qp12_d4;
    always @(posedge clk)
        n1008_q <= qp12_d5;
    always @(posedge clk)
        n1009_q <= qp12_d6;
    always @(posedge clk)
        n1010_q <= qp12_d7;
    always @(posedge clk)
        n1011_q <= qp12_d8;
    always @(posedge clk)
        n1012_q <= qm12;
    always @(posedge clk)
        n1013_q <= qm12_d1;
    always @(posedge clk)
        n1014_q <= qm12_d2;
    always @(posedge clk)
        n1015_q <= qm12_d3;
    always @(posedge clk)
        n1016_q <= qm12_d4;
    always @(posedge clk)
        n1017_q <= qm12_d5;
    always @(posedge clk)
        n1018_q <= qm12_d6;
    always @(posedge clk)
        n1019_q <= qm12_d7;
    always @(posedge clk)
        n1020_q <= qm12_d8;
    always @(posedge clk)
        n1021_q <= qm12_d9;
    always @(posedge clk)
        n1022_q <= qp11;
    always @(posedge clk)
        n1023_q <= qp11_d1;
    always @(posedge clk)
        n1024_q <= qp11_d2;
    always @(posedge clk)
        n1025_q <= qp11_d3;
    always @(posedge clk)
        n1026_q <= qp11_d4;
    always @(posedge clk)
        n1027_q <= qp11_d5;
    always @(posedge clk)
        n1028_q <= qp11_d6;
    always @(posedge clk)
        n1029_q <= qp11_d7;
    always @(posedge clk)
        n1030_q <= qm11;
    always @(posedge clk)
        n1031_q <= qm11_d1;
    always @(posedge clk)
        n1032_q <= qm11_d2;
    always @(posedge clk)
        n1033_q <= qm11_d3;
    always @(posedge clk)
        n1034_q <= qm11_d4;
    always @(posedge clk)
        n1035_q <= qm11_d5;
    always @(posedge clk)
        n1036_q <= qm11_d6;
    always @(posedge clk)
        n1037_q <= qm11_d7;
    always @(posedge clk)
        n1038_q <= qm11_d8;
    always @(posedge clk)
        n1039_q <= qp10;
    always @(posedge clk)
        n1040_q <= qp10_d1;
    always @(posedge clk)
        n1041_q <= qp10_d2;
    always @(posedge clk)
        n1042_q <= qp10_d3;
    always @(posedge clk)
        n1043_q <= qp10_d4;
    always @(posedge clk)
        n1044_q <= qp10_d5;
    always @(posedge clk)
        n1045_q <= qp10_d6;
    always @(posedge clk)
        n1046_q <= qp10_d7;
    always @(posedge clk)
        n1047_q <= qm10;
    always @(posedge clk)
        n1048_q <= qm10_d1;
    always @(posedge clk)
        n1049_q <= qm10_d2;
    always @(posedge clk)
        n1050_q <= qm10_d3;
    always @(posedge clk)
        n1051_q <= qm10_d4;
    always @(posedge clk)
        n1052_q <= qm10_d5;
    always @(posedge clk)
        n1053_q <= qm10_d6;
    always @(posedge clk)
        n1054_q <= qm10_d7;
    always @(posedge clk)
        n1055_q <= qm10_d8;
    always @(posedge clk)
        n1056_q <= qp9;
    always @(posedge clk)
        n1057_q <= qp9_d1;
    always @(posedge clk)
        n1058_q <= qp9_d2;
    always @(posedge clk)
        n1059_q <= qp9_d3;
    always @(posedge clk)
        n1060_q <= qp9_d4;
    always @(posedge clk)
        n1061_q <= qp9_d5;
    always @(posedge clk)
        n1062_q <= qp9_d6;
    always @(posedge clk)
        n1063_q <= qm9;
    always @(posedge clk)
        n1064_q <= qm9_d1;
    always @(posedge clk)
        n1065_q <= qm9_d2;
    always @(posedge clk)
        n1066_q <= qm9_d3;
    always @(posedge clk)
        n1067_q <= qm9_d4;
    always @(posedge clk)
        n1068_q <= qm9_d5;
    always @(posedge clk)
        n1069_q <= qm9_d6;
    always @(posedge clk)
        n1070_q <= qm9_d7;
    always @(posedge clk)
        n1071_q <= qp8;
    always @(posedge clk)
        n1072_q <= qp8_d1;
    always @(posedge clk)
        n1073_q <= qp8_d2;
    always @(posedge clk)
        n1074_q <= qp8_d3;
    always @(posedge clk)
        n1075_q <= qp8_d4;
    always @(posedge clk)
        n1076_q <= qp8_d5;
    always @(posedge clk)
        n1077_q <= qm8;
    always @(posedge clk)
        n1078_q <= qm8_d1;
    always @(posedge clk)
        n1079_q <= qm8_d2;
    always @(posedge clk)
        n1080_q <= qm8_d3;
    always @(posedge clk)
        n1081_q <= qm8_d4;
    always @(posedge clk)
        n1082_q <= qm8_d5;
    always @(posedge clk)
        n1083_q <= qm8_d6;
    always @(posedge clk)
        n1084_q <= qp7;
    always @(posedge clk)
        n1085_q <= qp7_d1;
    always @(posedge clk)
        n1086_q <= qp7_d2;
    always @(posedge clk)
        n1087_q <= qp7_d3;
    always @(posedge clk)
        n1088_q <= qp7_d4;
    always @(posedge clk)
        n1089_q <= qm7;
    always @(posedge clk)
        n1090_q <= qm7_d1;
    always @(posedge clk)
        n1091_q <= qm7_d2;
    always @(posedge clk)
        n1092_q <= qm7_d3;
    always @(posedge clk)
        n1093_q <= qm7_d4;
    always @(posedge clk)
        n1094_q <= qm7_d5;
    always @(posedge clk)
        n1095_q <= qp6;
    always @(posedge clk)
        n1096_q <= qp6_d1;
    always @(posedge clk)
        n1097_q <= qp6_d2;
    always @(posedge clk)
        n1098_q <= qp6_d3;
    always @(posedge clk)
        n1099_q <= qm6;
    always @(posedge clk)
        n1100_q <= qm6_d1;
    always @(posedge clk)
        n1101_q <= qm6_d2;
    always @(posedge clk)
        n1102_q <= qm6_d3;
    always @(posedge clk)
        n1103_q <= qm6_d4;
    always @(posedge clk)
        n1104_q <= qp5;
    always @(posedge clk)
        n1105_q <= qp5_d1;
    always @(posedge clk)
        n1106_q <= qp5_d2;
    always @(posedge clk)
        n1107_q <= qm5;
    always @(posedge clk)
        n1108_q <= qm5_d1;
    always @(posedge clk)
        n1109_q <= qm5_d2;
    always @(posedge clk)
        n1110_q <= qm5_d3;
    always @(posedge clk)
        n1111_q <= qp4;
    always @(posedge clk)
        n1112_q <= qp4_d1;
    always @(posedge clk)
        n1113_q <= qm4;
    always @(posedge clk)
        n1114_q <= qm4_d1;
    always @(posedge clk)
        n1115_q <= qm4_d2;
    always @(posedge clk)
        n1116_q <= qp3;
    always @(posedge clk)
        n1117_q <= qm3;
    always @(posedge clk)
        n1118_q <= qm3_d1;
    always @(posedge clk)
        n1119_q <= qp2;
    always @(posedge clk)
        n1120_q <= qm2;
    always @(posedge clk)
        n1121_q <= qm2_d1;
    always @(posedge clk)
        n1122_q <= qm1;
    always @(posedge clk)
        n1123_q <= qp;
endmodule

