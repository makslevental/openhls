module fsqrt
  (input wire clk,
   input wire [18:0] X,
   output wire [18:0] R);
  wire [10:0] fracx;
  wire [4:0] ern0;
  wire [2:0] xsx;
  wire [4:0] ern1;
  wire [4:0] ern1_d1;
  wire [4:0] ern1_d2;
  wire [4:0] ern1_d3;
  wire [14:0] fracxnorm;
  wire [1:0] s0;
  wire [14:0] t1;
  wire d1;
  wire [15:0] t1s;
  wire [5:0] t1s_h;
  wire [9:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [14:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [15:0] t2s;
  wire [6:0] t2s_h;
  wire [8:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [14:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [15:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [7:0] t3s_l;
  wire [7:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [14:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [15:0] t4s;
  wire [8:0] t4s_h;
  wire [6:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [14:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [15:0] t5s;
  wire [9:0] t5s_h;
  wire [5:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [14:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [15:0] t6s;
  wire [10:0] t6s_h;
  wire [4:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [14:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [15:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire [3:0] t7s_l;
  wire [3:0] t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [14:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [15:0] t8s;
  wire [12:0] t8s_h;
  wire [2:0] t8s_l;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [14:0] t9;
  wire [9:0] s8;
  wire d9;
  wire [15:0] t9s;
  wire [13:0] t9s_h;
  wire [1:0] t9s_l;
  wire [13:0] u9;
  wire [13:0] t11_h;
  wire [14:0] t10;
  wire [10:0] s9;
  wire d10;
  wire d10_d1;
  wire [15:0] t10s;
  wire [14:0] t10s_h;
  wire [14:0] t10s_h_d1;
  wire t10s_l;
  wire t10s_l_d1;
  wire [14:0] u10;
  wire [14:0] u10_d1;
  wire [14:0] t12_h;
  wire [14:0] t11;
  wire [11:0] s10;
  wire [11:0] s10_d1;
  wire d11;
  wire [15:0] t11s;
  wire [15:0] t11s_h;
  wire [15:0] u11;
  wire [15:0] t13_h;
  wire [14:0] t12;
  wire [12:0] s11;
  wire d13;
  wire [13:0] mr;
  wire [10:0] fr;
  wire round;
  wire [10:0] frrnd;
  wire [15:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [2:0] xsr_d3;
  wire [10:0] n26_o;
  wire [3:0] n27_o;
  wire [4:0] n29_o;
  wire [2:0] n30_o;
  wire [4:0] n32_o;
  wire n33_o;
  wire [4:0] n34_o;
  wire [4:0] n35_o;
  wire [11:0] n37_o;
  wire [14:0] n39_o;
  wire n40_o;
  wire n41_o;
  wire [14:0] n42_o;
  wire [12:0] n44_o;
  wire [14:0] n46_o;
  wire [3:0] n48_o;
  wire [3:0] n50_o;
  wire [10:0] n51_o;
  wire [14:0] n52_o;
  wire n53_o;
  wire n54_o;
  wire [15:0] n56_o;
  wire [5:0] n57_o;
  wire [9:0] n58_o;
  wire [2:0] n60_o;
  wire [3:0] n61_o;
  wire n62_o;
  wire [4:0] n63_o;
  wire [5:0] n65_o;
  wire [5:0] n66_o;
  wire [5:0] n67_o;
  wire [5:0] n68_o;
  wire [4:0] n69_o;
  wire [14:0] n70_o;
  wire [2:0] n71_o;
  wire n72_o;
  wire n73_o;
  wire [15:0] n75_o;
  wire [6:0] n76_o;
  wire [8:0] n77_o;
  wire [3:0] n79_o;
  wire [4:0] n80_o;
  wire n81_o;
  wire [5:0] n82_o;
  wire [6:0] n84_o;
  wire [6:0] n85_o;
  wire [6:0] n86_o;
  wire [6:0] n87_o;
  wire [5:0] n88_o;
  wire [14:0] n89_o;
  wire [3:0] n90_o;
  wire n91_o;
  wire n92_o;
  wire [15:0] n94_o;
  wire [7:0] n95_o;
  wire [7:0] n96_o;
  wire [4:0] n98_o;
  wire [5:0] n99_o;
  wire n100_o;
  wire [6:0] n101_o;
  wire [7:0] n103_o;
  wire [7:0] n104_o;
  wire [7:0] n105_o;
  wire [7:0] n106_o;
  wire [6:0] n107_o;
  wire [14:0] n108_o;
  wire [4:0] n109_o;
  wire n110_o;
  wire n111_o;
  wire [15:0] n113_o;
  wire [8:0] n114_o;
  wire [6:0] n115_o;
  wire [5:0] n117_o;
  wire [6:0] n118_o;
  wire n119_o;
  wire [7:0] n120_o;
  wire [8:0] n122_o;
  wire [8:0] n123_o;
  wire [8:0] n124_o;
  wire [8:0] n125_o;
  wire [7:0] n126_o;
  wire [14:0] n127_o;
  wire [5:0] n128_o;
  wire n129_o;
  wire n130_o;
  wire [15:0] n132_o;
  wire [9:0] n133_o;
  wire [5:0] n134_o;
  wire [6:0] n136_o;
  wire [7:0] n137_o;
  wire n138_o;
  wire [8:0] n139_o;
  wire [9:0] n141_o;
  wire [9:0] n142_o;
  wire [9:0] n143_o;
  wire [9:0] n144_o;
  wire [8:0] n145_o;
  wire [14:0] n146_o;
  wire [6:0] n147_o;
  wire n148_o;
  wire n149_o;
  wire [15:0] n151_o;
  wire [10:0] n152_o;
  wire [4:0] n153_o;
  wire [7:0] n155_o;
  wire [8:0] n156_o;
  wire n157_o;
  wire [9:0] n158_o;
  wire [10:0] n160_o;
  wire [10:0] n161_o;
  wire [10:0] n162_o;
  wire [10:0] n163_o;
  wire [9:0] n164_o;
  wire [14:0] n165_o;
  wire [7:0] n166_o;
  wire n167_o;
  wire n168_o;
  wire [15:0] n170_o;
  wire [11:0] n171_o;
  wire [3:0] n172_o;
  wire [8:0] n174_o;
  wire [9:0] n175_o;
  wire n176_o;
  wire [10:0] n177_o;
  wire [11:0] n179_o;
  wire [11:0] n180_o;
  wire [11:0] n181_o;
  wire [11:0] n182_o;
  wire [10:0] n183_o;
  wire [14:0] n184_o;
  wire [8:0] n185_o;
  wire n186_o;
  wire n187_o;
  wire [15:0] n189_o;
  wire [12:0] n190_o;
  wire [2:0] n191_o;
  wire [9:0] n193_o;
  wire [10:0] n194_o;
  wire n195_o;
  wire [11:0] n196_o;
  wire [12:0] n198_o;
  wire [12:0] n199_o;
  wire [12:0] n200_o;
  wire [12:0] n201_o;
  wire [11:0] n202_o;
  wire [14:0] n203_o;
  wire [9:0] n204_o;
  wire n205_o;
  wire n206_o;
  wire [15:0] n208_o;
  wire [13:0] n209_o;
  wire [1:0] n210_o;
  wire [10:0] n212_o;
  wire [11:0] n213_o;
  wire n214_o;
  wire [12:0] n215_o;
  wire [13:0] n217_o;
  wire [13:0] n218_o;
  wire [13:0] n219_o;
  wire [13:0] n220_o;
  wire [12:0] n221_o;
  wire [14:0] n222_o;
  wire [10:0] n223_o;
  wire n224_o;
  wire n225_o;
  wire [15:0] n227_o;
  wire [14:0] n228_o;
  wire n229_o;
  wire [11:0] n231_o;
  wire [12:0] n232_o;
  wire n233_o;
  wire [13:0] n234_o;
  wire [14:0] n236_o;
  wire [14:0] n237_o;
  wire [14:0] n238_o;
  wire [14:0] n239_o;
  wire [13:0] n240_o;
  wire [14:0] n241_o;
  wire [11:0] n242_o;
  wire n243_o;
  wire n244_o;
  wire [15:0] n246_o;
  wire [12:0] n248_o;
  wire [13:0] n249_o;
  wire n250_o;
  wire [14:0] n251_o;
  wire [15:0] n253_o;
  wire [15:0] n254_o;
  wire [15:0] n255_o;
  wire [15:0] n256_o;
  wire [14:0] n257_o;
  wire [12:0] n258_o;
  wire n259_o;
  wire n260_o;
  wire [13:0] n261_o;
  wire [10:0] n262_o;
  wire n263_o;
  wire [10:0] n265_o;
  wire [10:0] n266_o;
  wire [15:0] n267_o;
  wire n270_o;
  wire n273_o;
  wire n276_o;
  wire n279_o;
  wire [3:0] n281_o;
  reg [2:0] n282_o;
  wire [18:0] n283_o;
  reg [4:0] n284_q;
  reg [4:0] n285_q;
  reg [4:0] n286_q;
  reg n287_q;
  reg [7:0] n288_q;
  reg [7:0] n289_q;
  reg [7:0] n290_q;
  reg [4:0] n291_q;
  reg n292_q;
  reg [11:0] n293_q;
  reg [3:0] n294_q;
  reg [11:0] n295_q;
  reg [8:0] n296_q;
  reg n297_q;
  reg [14:0] n298_q;
  reg n299_q;
  reg [14:0] n300_q;
  reg [11:0] n301_q;
  reg [2:0] n302_q;
  reg [2:0] n303_q;
  reg [2:0] n304_q;
  assign R = n283_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:30:8  */
  assign fracx = n26_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:31:8  */
  assign ern0 = n29_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:32:8  */
  assign xsx = n30_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:33:8  */
  assign ern1 = n35_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:33:14  */
  assign ern1_d1 = n284_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:33:23  */
  assign ern1_d2 = n285_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:33:32  */
  assign ern1_d3 = n286_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:34:8  */
  assign fracxnorm = n42_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:36:8  */
  assign t1 = n52_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:37:8  */
  assign d1 = n54_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:38:8  */
  assign t1s = n56_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:39:8  */
  assign t1s_h = n57_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:40:8  */
  assign t1s_l = n58_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:41:8  */
  assign u1 = n65_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:42:8  */
  assign t3_h = n67_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:43:8  */
  assign t2 = n70_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:44:8  */
  assign s1 = n71_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:45:8  */
  assign d2 = n73_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:46:8  */
  assign t2s = n75_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:47:8  */
  assign t2s_h = n76_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:48:8  */
  assign t2s_l = n77_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:49:8  */
  assign u2 = n84_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:50:8  */
  assign t4_h = n86_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:51:8  */
  assign t3 = n89_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:52:8  */
  assign s2 = n90_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:53:8  */
  assign d3 = n92_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:53:12  */
  assign d3_d1 = n287_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:54:8  */
  assign t3s = n94_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:55:8  */
  assign t3s_h = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:55:15  */
  assign t3s_h_d1 = n288_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:56:8  */
  assign t3s_l = n96_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:56:15  */
  assign t3s_l_d1 = n289_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:57:8  */
  assign u3 = n103_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:57:12  */
  assign u3_d1 = n290_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:58:8  */
  assign t5_h = n105_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:59:8  */
  assign t4 = n108_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:60:8  */
  assign s3 = n109_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:60:12  */
  assign s3_d1 = n291_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:61:8  */
  assign d4 = n111_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:62:8  */
  assign t4s = n113_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:63:8  */
  assign t4s_h = n114_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:64:8  */
  assign t4s_l = n115_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:65:8  */
  assign u4 = n122_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:66:8  */
  assign t6_h = n124_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:67:8  */
  assign t5 = n127_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:68:8  */
  assign s4 = n128_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:69:8  */
  assign d5 = n130_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:70:8  */
  assign t5s = n132_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:71:8  */
  assign t5s_h = n133_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:72:8  */
  assign t5s_l = n134_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:73:8  */
  assign u5 = n141_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:74:8  */
  assign t7_h = n143_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:75:8  */
  assign t6 = n146_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:76:8  */
  assign s5 = n147_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:77:8  */
  assign d6 = n149_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:78:8  */
  assign t6s = n151_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:79:8  */
  assign t6s_h = n152_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:80:8  */
  assign t6s_l = n153_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:81:8  */
  assign u6 = n160_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:82:8  */
  assign t8_h = n162_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:83:8  */
  assign t7 = n165_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:84:8  */
  assign s6 = n166_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:85:8  */
  assign d7 = n168_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:85:12  */
  assign d7_d1 = n292_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:86:8  */
  assign t7s = n170_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:87:8  */
  assign t7s_h = n171_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:87:15  */
  assign t7s_h_d1 = n293_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:88:8  */
  assign t7s_l = n172_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:88:15  */
  assign t7s_l_d1 = n294_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:89:8  */
  assign u7 = n179_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:89:12  */
  assign u7_d1 = n295_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:90:8  */
  assign t9_h = n181_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:91:8  */
  assign t8 = n184_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:92:8  */
  assign s7 = n185_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:92:12  */
  assign s7_d1 = n296_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:93:8  */
  assign d8 = n187_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:94:8  */
  assign t8s = n189_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:95:8  */
  assign t8s_h = n190_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:96:8  */
  assign t8s_l = n191_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:97:8  */
  assign u8 = n198_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:98:8  */
  assign t10_h = n200_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:99:8  */
  assign t9 = n203_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:100:8  */
  assign s8 = n204_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:101:8  */
  assign d9 = n206_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:102:8  */
  assign t9s = n208_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:103:8  */
  assign t9s_h = n209_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:104:8  */
  assign t9s_l = n210_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:105:8  */
  assign u9 = n217_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:106:8  */
  assign t11_h = n219_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:107:8  */
  assign t10 = n222_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:108:8  */
  assign s9 = n223_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:109:8  */
  assign d10 = n225_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:109:13  */
  assign d10_d1 = n297_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:110:8  */
  assign t10s = n227_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:111:8  */
  assign t10s_h = n228_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:111:16  */
  assign t10s_h_d1 = n298_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:112:8  */
  assign t10s_l = n229_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:112:16  */
  assign t10s_l_d1 = n299_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:113:8  */
  assign u10 = n236_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:113:13  */
  assign u10_d1 = n300_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:114:8  */
  assign t12_h = n238_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:115:8  */
  assign t11 = n241_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:116:8  */
  assign s10 = n242_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:116:13  */
  assign s10_d1 = n301_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:117:8  */
  assign d11 = n244_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:271:18  */
  assign t11s = n246_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:119:8  */
  assign t11s_h = t11s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:120:8  */
  assign u11 = n253_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:121:8  */
  assign t13_h = n255_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:122:8  */
  assign t12 = n257_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:123:8  */
  assign s11 = n258_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:124:8  */
  assign d13 = n260_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:125:8  */
  assign mr = n261_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:126:8  */
  assign fr = n262_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:127:8  */
  assign round = n263_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:128:8  */
  assign frrnd = n266_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:129:8  */
  assign rn2 = n267_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:130:8  */
  assign xsr = n282_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:130:13  */
  assign xsr_d1 = n302_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:130:21  */
  assign xsr_d2 = n303_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:130:29  */
  assign xsr_d3 = n304_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:158:14  */
  assign n26_o = X[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:159:19  */
  assign n27_o = X[15:12];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:159:16  */
  assign n29_o = {1'b0, n27_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:160:12  */
  assign n30_o = X[18:16];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:161:17  */
  assign n32_o = ern0 + 5'b00111;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:161:51  */
  assign n33_o = X[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:161:48  */
  assign n34_o = {4'b0, n33_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:161:48  */
  assign n35_o = n32_o + n34_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:162:21  */
  assign n37_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:162:29  */
  assign n39_o = {n37_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:162:43  */
  assign n40_o = X[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:162:48  */
  assign n41_o = ~n40_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:162:37  */
  assign n42_o = n41_o ? n39_o : n46_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:163:15  */
  assign n44_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:163:22  */
  assign n46_o = {n44_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:165:29  */
  assign n48_o = fracxnorm[14:11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:165:18  */
  assign n50_o = 4'b0111 + n48_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:165:56  */
  assign n51_o = fracxnorm[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:165:45  */
  assign n52_o = {n50_o, n51_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:169:16  */
  assign n53_o = t1[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:169:10  */
  assign n54_o = ~n53_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:170:14  */
  assign n56_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:171:16  */
  assign n57_o = t1s[15:10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:172:16  */
  assign n58_o = t1s[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:173:15  */
  assign n60_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:173:20  */
  assign n61_o = {n60_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:173:28  */
  assign n62_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:173:25  */
  assign n63_o = {n61_o, n62_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:173:36  */
  assign n65_o = {n63_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:174:20  */
  assign n66_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:174:25  */
  assign n67_o = d1 ? n66_o : n68_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:175:20  */
  assign n68_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:176:14  */
  assign n69_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:176:27  */
  assign n70_o = {n69_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:177:13  */
  assign n71_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:179:16  */
  assign n72_o = t2[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:179:10  */
  assign n73_o = ~n72_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:180:14  */
  assign n75_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:181:16  */
  assign n76_o = t2s[15:9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:182:16  */
  assign n77_o = t2s[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:183:15  */
  assign n79_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:183:20  */
  assign n80_o = {n79_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:183:28  */
  assign n81_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:183:25  */
  assign n82_o = {n80_o, n81_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:183:36  */
  assign n84_o = {n82_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:184:20  */
  assign n85_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:184:25  */
  assign n86_o = d2 ? n85_o : n87_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:185:20  */
  assign n87_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:186:14  */
  assign n88_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:186:27  */
  assign n89_o = {n88_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:187:13  */
  assign n90_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:189:16  */
  assign n91_o = t3[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:189:10  */
  assign n92_o = ~n91_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:190:14  */
  assign n94_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:191:16  */
  assign n95_o = t3s[15:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:192:16  */
  assign n96_o = t3s[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:193:15  */
  assign n98_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:193:20  */
  assign n99_o = {n98_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:193:28  */
  assign n100_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:193:25  */
  assign n101_o = {n99_o, n100_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:193:36  */
  assign n103_o = {n101_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:194:23  */
  assign n104_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:194:31  */
  assign n105_o = d3_d1 ? n104_o : n106_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:195:23  */
  assign n106_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:196:14  */
  assign n107_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:196:27  */
  assign n108_o = {n107_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:197:13  */
  assign n109_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:199:16  */
  assign n110_o = t4[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:199:10  */
  assign n111_o = ~n110_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:200:14  */
  assign n113_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:201:16  */
  assign n114_o = t4s[15:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:202:16  */
  assign n115_o = t4s[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:203:15  */
  assign n117_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:203:23  */
  assign n118_o = {n117_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:203:31  */
  assign n119_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:203:28  */
  assign n120_o = {n118_o, n119_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:203:39  */
  assign n122_o = {n120_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:204:20  */
  assign n123_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:204:25  */
  assign n124_o = d4 ? n123_o : n125_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:205:20  */
  assign n125_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:206:14  */
  assign n126_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:206:27  */
  assign n127_o = {n126_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:207:16  */
  assign n128_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:209:16  */
  assign n129_o = t5[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:209:10  */
  assign n130_o = ~n129_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:210:14  */
  assign n132_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:211:16  */
  assign n133_o = t5s[15:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:212:16  */
  assign n134_o = t5s[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:213:15  */
  assign n136_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:213:20  */
  assign n137_o = {n136_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:213:28  */
  assign n138_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:213:25  */
  assign n139_o = {n137_o, n138_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:213:36  */
  assign n141_o = {n139_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:214:20  */
  assign n142_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:214:25  */
  assign n143_o = d5 ? n142_o : n144_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:215:20  */
  assign n144_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:216:14  */
  assign n145_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:216:27  */
  assign n146_o = {n145_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:217:13  */
  assign n147_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:219:16  */
  assign n148_o = t6[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:219:10  */
  assign n149_o = ~n148_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:220:14  */
  assign n151_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:221:16  */
  assign n152_o = t6s[15:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:222:16  */
  assign n153_o = t6s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:223:15  */
  assign n155_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:223:20  */
  assign n156_o = {n155_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:223:28  */
  assign n157_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:223:25  */
  assign n158_o = {n156_o, n157_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:223:36  */
  assign n160_o = {n158_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:224:20  */
  assign n161_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:224:25  */
  assign n162_o = d6 ? n161_o : n163_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:225:20  */
  assign n163_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:226:14  */
  assign n164_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:226:27  */
  assign n165_o = {n164_o, t6s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:227:13  */
  assign n166_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:229:16  */
  assign n167_o = t7[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:229:10  */
  assign n168_o = ~n167_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:230:14  */
  assign n170_o = {t7, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:231:16  */
  assign n171_o = t7s[15:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:232:16  */
  assign n172_o = t7s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:233:15  */
  assign n174_o = {1'b0, s6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:233:20  */
  assign n175_o = {n174_o, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:233:28  */
  assign n176_o = ~d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:233:25  */
  assign n177_o = {n175_o, n176_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:233:36  */
  assign n179_o = {n177_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:234:23  */
  assign n180_o = t7s_h_d1 - u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:234:31  */
  assign n181_o = d7_d1 ? n180_o : n182_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:235:23  */
  assign n182_o = t7s_h_d1 + u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:236:14  */
  assign n183_o = t9_h[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:236:28  */
  assign n184_o = {n183_o, t7s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:237:13  */
  assign n185_o = {s6, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:239:16  */
  assign n186_o = t8[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:239:10  */
  assign n187_o = ~n186_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:240:14  */
  assign n189_o = {t8, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:241:16  */
  assign n190_o = t8s[15:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:242:16  */
  assign n191_o = t8s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:243:15  */
  assign n193_o = {1'b0, s7_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:243:23  */
  assign n194_o = {n193_o, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:243:31  */
  assign n195_o = ~d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:243:28  */
  assign n196_o = {n194_o, n195_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:243:39  */
  assign n198_o = {n196_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:244:21  */
  assign n199_o = t8s_h - u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:244:26  */
  assign n200_o = d8 ? n199_o : n201_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:245:20  */
  assign n201_o = t8s_h + u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:246:15  */
  assign n202_o = t10_h[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:246:29  */
  assign n203_o = {n202_o, t8s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:247:16  */
  assign n204_o = {s7_d1, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:249:16  */
  assign n205_o = t9[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:249:10  */
  assign n206_o = ~n205_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:250:14  */
  assign n208_o = {t9, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:251:16  */
  assign n209_o = t9s[15:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:252:16  */
  assign n210_o = t9s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:253:15  */
  assign n212_o = {1'b0, s8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:253:20  */
  assign n213_o = {n212_o, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:253:28  */
  assign n214_o = ~d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:253:25  */
  assign n215_o = {n213_o, n214_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:253:36  */
  assign n217_o = {n215_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:254:21  */
  assign n218_o = t9s_h - u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:254:26  */
  assign n219_o = d9 ? n218_o : n220_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:255:20  */
  assign n220_o = t9s_h + u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:256:16  */
  assign n221_o = t11_h[12:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:256:30  */
  assign n222_o = {n221_o, t9s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:257:13  */
  assign n223_o = {s8, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:259:18  */
  assign n224_o = t10[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:259:11  */
  assign n225_o = ~n224_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:260:16  */
  assign n227_o = {t10, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:261:18  */
  assign n228_o = t10s[15:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:262:18  */
  assign n229_o = t10s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:263:16  */
  assign n231_o = {1'b0, s9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:263:21  */
  assign n232_o = {n231_o, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:263:30  */
  assign n233_o = ~d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:263:27  */
  assign n234_o = {n232_o, n233_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:263:39  */
  assign n236_o = {n234_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:264:25  */
  assign n237_o = t10s_h_d1 - u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:264:34  */
  assign n238_o = d10_d1 ? n237_o : n239_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:265:24  */
  assign n239_o = t10s_h_d1 + u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:266:16  */
  assign n240_o = t12_h[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:266:30  */
  assign n241_o = {n240_o, t10s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:267:14  */
  assign n242_o = {s9, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:269:18  */
  assign n243_o = t11[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:269:11  */
  assign n244_o = ~n243_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:270:16  */
  assign n246_o = {t11, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:272:16  */
  assign n248_o = {1'b0, s10_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:272:25  */
  assign n249_o = {n248_o, d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:272:34  */
  assign n250_o = ~d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:272:31  */
  assign n251_o = {n249_o, n250_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:272:43  */
  assign n253_o = {n251_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:273:22  */
  assign n254_o = t11s_h - u11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:273:28  */
  assign n255_o = d11 ? n254_o : n256_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:274:21  */
  assign n256_o = t11s_h + u11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:275:16  */
  assign n257_o = t13_h[14:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:276:18  */
  assign n258_o = {s10_d1, d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:277:18  */
  assign n259_o = t12[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:277:11  */
  assign n260_o = ~n259_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:278:14  */
  assign n261_o = {s11, d13};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:279:12  */
  assign n262_o = mr[11:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:280:15  */
  assign n263_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:281:40  */
  assign n265_o = {10'b0000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:281:16  */
  assign n266_o = fr + n265_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:282:19  */
  assign n267_o = {ern1_d3, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:285:21  */
  assign n270_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:286:21  */
  assign n273_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:287:21  */
  assign n276_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:288:21  */
  assign n279_o = xsx == 3'b001;
  assign n281_o = {n279_o, n276_o, n273_o, n270_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:284:4  */
  always @*
    case (n281_o)
      4'b1000: n282_o = 3'b001;
      4'b0100: n282_o = 3'b000;
      4'b0010: n282_o = 3'b100;
      4'b0001: n282_o = 3'b010;
      default: n282_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:290:16  */
  assign n283_o = {xsr_d3, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n284_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n285_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n286_q <= ern1_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n287_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n288_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n289_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n290_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n291_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n292_q <= d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n293_q <= t7s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n294_q <= t7s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n295_q <= u7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n296_q <= s7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n297_q <= d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n298_q <= t10s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n299_q <= t10s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n300_q <= u10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n301_q <= s10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n302_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n303_q <= xsr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_5_11.vhdl:134:10  */
  always @(posedge clk)
    n304_q <= xsr_d2;
endmodule

