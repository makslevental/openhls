module fsqrt#(parameter ID=1)
  (input  clk,
   input  [18:0] X,
   output [18:0] R);
  wire [7:0] fracx;
  wire [7:0] ern0;
  wire [2:0] xsx;
  wire [7:0] ern1;
  wire [7:0] ern1_d1;
  wire [7:0] ern1_d2;
  wire [11:0] fracxnorm;
  wire [1:0] s0;
  wire [11:0] t1;
  wire d1;
  wire [12:0] t1s;
  wire [5:0] t1s_h;
  wire [6:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [11:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [12:0] t2s;
  wire [6:0] t2s_h;
  wire [5:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [11:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [12:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [4:0] t3s_l;
  wire [4:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [11:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [12:0] t4s;
  wire [8:0] t4s_h;
  wire [3:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [11:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [12:0] t5s;
  wire [9:0] t5s_h;
  wire [2:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [11:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [12:0] t6s;
  wire [10:0] t6s_h;
  wire [1:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [11:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [12:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire t7s_l;
  wire t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [11:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [12:0] t8s;
  wire [12:0] t8s_h;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [11:0] t9;
  wire [9:0] s8;
  wire d10;
  wire [10:0] mr;
  wire [7:0] fr;
  wire round;
  wire [7:0] frrnd;
  wire [15:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [7:0] n19_o;
  wire [6:0] n20_o;
  wire [7:0] n22_o;
  wire [2:0] n23_o;
  wire [7:0] n25_o;
  wire n26_o;
  wire [7:0] n27_o;
  wire [7:0] n28_o;
  wire [8:0] n30_o;
  wire [11:0] n32_o;
  wire n33_o;
  wire n34_o;
  wire [11:0] n35_o;
  wire [9:0] n37_o;
  wire [11:0] n39_o;
  wire [3:0] n41_o;
  wire [3:0] n43_o;
  wire [7:0] n44_o;
  wire [11:0] n45_o;
  wire n46_o;
  wire n47_o;
  wire [12:0] n49_o;
  wire [5:0] n50_o;
  wire [6:0] n51_o;
  wire [2:0] n53_o;
  wire [3:0] n54_o;
  wire n55_o;
  wire [4:0] n56_o;
  wire [5:0] n58_o;
  wire [5:0] n59_o;
  wire [5:0] n60_o;
  wire [5:0] n61_o;
  wire [4:0] n62_o;
  wire [11:0] n63_o;
  wire [2:0] n64_o;
  wire n65_o;
  wire n66_o;
  wire [12:0] n68_o;
  wire [6:0] n69_o;
  wire [5:0] n70_o;
  wire [3:0] n72_o;
  wire [4:0] n73_o;
  wire n74_o;
  wire [5:0] n75_o;
  wire [6:0] n77_o;
  wire [6:0] n78_o;
  wire [6:0] n79_o;
  wire [6:0] n80_o;
  wire [5:0] n81_o;
  wire [11:0] n82_o;
  wire [3:0] n83_o;
  wire n84_o;
  wire n85_o;
  wire [12:0] n87_o;
  wire [7:0] n88_o;
  wire [4:0] n89_o;
  wire [4:0] n91_o;
  wire [5:0] n92_o;
  wire n93_o;
  wire [6:0] n94_o;
  wire [7:0] n96_o;
  wire [7:0] n97_o;
  wire [7:0] n98_o;
  wire [7:0] n99_o;
  wire [6:0] n100_o;
  wire [11:0] n101_o;
  wire [4:0] n102_o;
  wire n103_o;
  wire n104_o;
  wire [12:0] n106_o;
  wire [8:0] n107_o;
  wire [3:0] n108_o;
  wire [5:0] n110_o;
  wire [6:0] n111_o;
  wire n112_o;
  wire [7:0] n113_o;
  wire [8:0] n115_o;
  wire [8:0] n116_o;
  wire [8:0] n117_o;
  wire [8:0] n118_o;
  wire [7:0] n119_o;
  wire [11:0] n120_o;
  wire [5:0] n121_o;
  wire n122_o;
  wire n123_o;
  wire [12:0] n125_o;
  wire [9:0] n126_o;
  wire [2:0] n127_o;
  wire [6:0] n129_o;
  wire [7:0] n130_o;
  wire n131_o;
  wire [8:0] n132_o;
  wire [9:0] n134_o;
  wire [9:0] n135_o;
  wire [9:0] n136_o;
  wire [9:0] n137_o;
  wire [8:0] n138_o;
  wire [11:0] n139_o;
  wire [6:0] n140_o;
  wire n141_o;
  wire n142_o;
  wire [12:0] n144_o;
  wire [10:0] n145_o;
  wire [1:0] n146_o;
  wire [7:0] n148_o;
  wire [8:0] n149_o;
  wire n150_o;
  wire [9:0] n151_o;
  wire [10:0] n153_o;
  wire [10:0] n154_o;
  wire [10:0] n155_o;
  wire [10:0] n156_o;
  wire [9:0] n157_o;
  wire [11:0] n158_o;
  wire [7:0] n159_o;
  wire n160_o;
  wire n161_o;
  wire [12:0] n163_o;
  wire [11:0] n164_o;
  wire n165_o;
  wire [8:0] n167_o;
  wire [9:0] n168_o;
  wire n169_o;
  wire [10:0] n170_o;
  wire [11:0] n172_o;
  wire [11:0] n173_o;
  wire [11:0] n174_o;
  wire [11:0] n175_o;
  wire [10:0] n176_o;
  wire [11:0] n177_o;
  wire [8:0] n178_o;
  wire n179_o;
  wire n180_o;
  wire [12:0] n182_o;
  wire [9:0] n184_o;
  wire [10:0] n185_o;
  wire n186_o;
  wire [11:0] n187_o;
  wire [12:0] n189_o;
  wire [12:0] n190_o;
  wire [12:0] n191_o;
  wire [12:0] n192_o;
  wire [11:0] n193_o;
  wire [9:0] n194_o;
  wire n195_o;
  wire n196_o;
  wire [10:0] n197_o;
  wire [7:0] n198_o;
  wire n199_o;
  wire [7:0] n201_o;
  wire [7:0] n202_o;
  wire [15:0] n203_o;
  wire n206_o;
  wire n209_o;
  wire n212_o;
  wire n215_o;
  wire [3:0] n217_o;
  reg [2:0] n218_o;
  wire [18:0] n219_o;
  reg [7:0] n220_q;
  reg [7:0] n221_q;
  reg n222_q;
  reg [7:0] n223_q;
  reg [4:0] n224_q;
  reg [7:0] n225_q;
  reg [4:0] n226_q;
  reg n227_q;
  reg [11:0] n228_q;
  reg n229_q;
  reg [11:0] n230_q;
  reg [8:0] n231_q;
  reg [2:0] n232_q;
  reg [2:0] n233_q;
  assign R = n219_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:30:8  */
  assign fracx = n19_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:31:8  */
  assign ern0 = n22_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:32:8  */
  assign xsx = n23_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:33:8  */
  assign ern1 = n28_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:33:14  */
  assign ern1_d1 = n220_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:33:23  */
  assign ern1_d2 = n221_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:34:8  */
  assign fracxnorm = n35_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:36:8  */
  assign t1 = n45_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:37:8  */
  assign d1 = n47_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:38:8  */
  assign t1s = n49_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:39:8  */
  assign t1s_h = n50_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:40:8  */
  assign t1s_l = n51_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:41:8  */
  assign u1 = n58_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:42:8  */
  assign t3_h = n60_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:43:8  */
  assign t2 = n63_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:44:8  */
  assign s1 = n64_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:45:8  */
  assign d2 = n66_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:46:8  */
  assign t2s = n68_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:47:8  */
  assign t2s_h = n69_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:48:8  */
  assign t2s_l = n70_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:49:8  */
  assign u2 = n77_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:50:8  */
  assign t4_h = n79_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:51:8  */
  assign t3 = n82_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:52:8  */
  assign s2 = n83_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:53:8  */
  assign d3 = n85_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:53:12  */
  assign d3_d1 = n222_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:54:8  */
  assign t3s = n87_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:55:8  */
  assign t3s_h = n88_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:55:15  */
  assign t3s_h_d1 = n223_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:56:8  */
  assign t3s_l = n89_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:56:15  */
  assign t3s_l_d1 = n224_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:57:8  */
  assign u3 = n96_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:57:12  */
  assign u3_d1 = n225_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:58:8  */
  assign t5_h = n98_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:59:8  */
  assign t4 = n101_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:60:8  */
  assign s3 = n102_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:60:12  */
  assign s3_d1 = n226_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:61:8  */
  assign d4 = n104_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:62:8  */
  assign t4s = n106_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:63:8  */
  assign t4s_h = n107_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:64:8  */
  assign t4s_l = n108_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:65:8  */
  assign u4 = n115_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:66:8  */
  assign t6_h = n117_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:67:8  */
  assign t5 = n120_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:68:8  */
  assign s4 = n121_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:69:8  */
  assign d5 = n123_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:70:8  */
  assign t5s = n125_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:71:8  */
  assign t5s_h = n126_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:72:8  */
  assign t5s_l = n127_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:73:8  */
  assign u5 = n134_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:74:8  */
  assign t7_h = n136_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:75:8  */
  assign t6 = n139_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:76:8  */
  assign s5 = n140_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:77:8  */
  assign d6 = n142_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:78:8  */
  assign t6s = n144_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:79:8  */
  assign t6s_h = n145_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:80:8  */
  assign t6s_l = n146_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:81:8  */
  assign u6 = n153_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:82:8  */
  assign t8_h = n155_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:83:8  */
  assign t7 = n158_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:84:8  */
  assign s6 = n159_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:85:8  */
  assign d7 = n161_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:85:12  */
  assign d7_d1 = n227_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:86:8  */
  assign t7s = n163_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:87:8  */
  assign t7s_h = n164_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:87:15  */
  assign t7s_h_d1 = n228_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:88:8  */
  assign t7s_l = n165_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:88:15  */
  assign t7s_l_d1 = n229_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:89:8  */
  assign u7 = n172_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:89:12  */
  assign u7_d1 = n230_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:90:8  */
  assign t9_h = n174_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:91:8  */
  assign t8 = n177_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:92:8  */
  assign s7 = n178_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:92:12  */
  assign s7_d1 = n231_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:93:8  */
  assign d8 = n180_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:210:16  */
  assign t8s = n182_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:95:8  */
  assign t8s_h = t8s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:96:8  */
  assign u8 = n189_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:97:8  */
  assign t10_h = n191_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:98:8  */
  assign t9 = n193_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:99:8  */
  assign s8 = n194_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:100:8  */
  assign d10 = n196_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:101:8  */
  assign mr = n197_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:102:8  */
  assign fr = n198_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:103:8  */
  assign round = n199_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:104:8  */
  assign frrnd = n202_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:105:8  */
  assign rn2 = n203_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:106:8  */
  assign xsr = n218_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:106:13  */
  assign xsr_d1 = n232_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:106:21  */
  assign xsr_d2 = n233_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:127:14  */
  assign n19_o = X[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:128:19  */
  assign n20_o = X[15:9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:128:16  */
  assign n22_o = {1'b0, n20_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:129:12  */
  assign n23_o = X[18:16];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:130:17  */
  assign n25_o = ern0 + 8'b00111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:130:51  */
  assign n26_o = X[8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:130:48  */
  assign n27_o = {7'b0, n26_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:130:48  */
  assign n28_o = n25_o + n27_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:131:21  */
  assign n30_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:131:29  */
  assign n32_o = {n30_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:131:43  */
  assign n33_o = X[8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:131:47  */
  assign n34_o = ~n33_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:131:37  */
  assign n35_o = n34_o ? n32_o : n39_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:132:15  */
  assign n37_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:132:22  */
  assign n39_o = {n37_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:134:29  */
  assign n41_o = fracxnorm[11:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:134:18  */
  assign n43_o = 4'b0111 + n41_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:134:55  */
  assign n44_o = fracxnorm[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:134:44  */
  assign n45_o = {n43_o, n44_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:138:16  */
  assign n46_o = t1[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:138:10  */
  assign n47_o = ~n46_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:139:14  */
  assign n49_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:140:16  */
  assign n50_o = t1s[12:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:141:16  */
  assign n51_o = t1s[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:142:15  */
  assign n53_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:142:20  */
  assign n54_o = {n53_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:142:28  */
  assign n55_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:142:25  */
  assign n56_o = {n54_o, n55_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:142:36  */
  assign n58_o = {n56_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:143:20  */
  assign n59_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:143:25  */
  assign n60_o = d1 ? n59_o : n61_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:144:20  */
  assign n61_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:145:14  */
  assign n62_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:145:27  */
  assign n63_o = {n62_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:146:13  */
  assign n64_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:148:16  */
  assign n65_o = t2[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:148:10  */
  assign n66_o = ~n65_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:149:14  */
  assign n68_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:150:16  */
  assign n69_o = t2s[12:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:151:16  */
  assign n70_o = t2s[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:152:15  */
  assign n72_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:152:20  */
  assign n73_o = {n72_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:152:28  */
  assign n74_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:152:25  */
  assign n75_o = {n73_o, n74_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:152:36  */
  assign n77_o = {n75_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:153:20  */
  assign n78_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:153:25  */
  assign n79_o = d2 ? n78_o : n80_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:154:20  */
  assign n80_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:155:14  */
  assign n81_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:155:27  */
  assign n82_o = {n81_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:156:13  */
  assign n83_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:158:16  */
  assign n84_o = t3[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:158:10  */
  assign n85_o = ~n84_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:159:14  */
  assign n87_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:160:16  */
  assign n88_o = t3s[12:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:161:16  */
  assign n89_o = t3s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:162:15  */
  assign n91_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:162:20  */
  assign n92_o = {n91_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:162:28  */
  assign n93_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:162:25  */
  assign n94_o = {n92_o, n93_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:162:36  */
  assign n96_o = {n94_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:163:23  */
  assign n97_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:163:31  */
  assign n98_o = d3_d1 ? n97_o : n99_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:164:23  */
  assign n99_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:165:14  */
  assign n100_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:165:27  */
  assign n101_o = {n100_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:166:13  */
  assign n102_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:168:16  */
  assign n103_o = t4[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:168:10  */
  assign n104_o = ~n103_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:169:14  */
  assign n106_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:170:16  */
  assign n107_o = t4s[12:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:171:16  */
  assign n108_o = t4s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:172:15  */
  assign n110_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:172:23  */
  assign n111_o = {n110_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:172:31  */
  assign n112_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:172:28  */
  assign n113_o = {n111_o, n112_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:172:39  */
  assign n115_o = {n113_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:173:20  */
  assign n116_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:173:25  */
  assign n117_o = d4 ? n116_o : n118_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:174:20  */
  assign n118_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:175:14  */
  assign n119_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:175:27  */
  assign n120_o = {n119_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:176:16  */
  assign n121_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:178:16  */
  assign n122_o = t5[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:178:10  */
  assign n123_o = ~n122_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:179:14  */
  assign n125_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:180:16  */
  assign n126_o = t5s[12:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:181:16  */
  assign n127_o = t5s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:182:15  */
  assign n129_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:182:20  */
  assign n130_o = {n129_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:182:28  */
  assign n131_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:182:25  */
  assign n132_o = {n130_o, n131_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:182:36  */
  assign n134_o = {n132_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:183:20  */
  assign n135_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:183:25  */
  assign n136_o = d5 ? n135_o : n137_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:184:20  */
  assign n137_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:185:14  */
  assign n138_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:185:27  */
  assign n139_o = {n138_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:186:13  */
  assign n140_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:188:16  */
  assign n141_o = t6[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:188:10  */
  assign n142_o = ~n141_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:189:14  */
  assign n144_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:190:16  */
  assign n145_o = t6s[12:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:191:16  */
  assign n146_o = t6s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:192:15  */
  assign n148_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:192:20  */
  assign n149_o = {n148_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:192:28  */
  assign n150_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:192:25  */
  assign n151_o = {n149_o, n150_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:192:36  */
  assign n153_o = {n151_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:193:20  */
  assign n154_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:193:25  */
  assign n155_o = d6 ? n154_o : n156_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:194:20  */
  assign n156_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:195:14  */
  assign n157_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:195:27  */
  assign n158_o = {n157_o, t6s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:196:13  */
  assign n159_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:198:16  */
  assign n160_o = t7[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:198:10  */
  assign n161_o = ~n160_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:199:14  */
  assign n163_o = {t7, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:200:16  */
  assign n164_o = t7s[12:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:201:16  */
  assign n165_o = t7s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:202:15  */
  assign n167_o = {1'b0, s6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:202:20  */
  assign n168_o = {n167_o, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:202:28  */
  assign n169_o = ~d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:202:25  */
  assign n170_o = {n168_o, n169_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:202:36  */
  assign n172_o = {n170_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:203:23  */
  assign n173_o = t7s_h_d1 - u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:203:31  */
  assign n174_o = d7_d1 ? n173_o : n175_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:204:23  */
  assign n175_o = t7s_h_d1 + u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:205:14  */
  assign n176_o = t9_h[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:205:28  */
  assign n177_o = {n176_o, t7s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:206:13  */
  assign n178_o = {s6, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:208:16  */
  assign n179_o = t8[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:208:10  */
  assign n180_o = ~n179_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:209:14  */
  assign n182_o = {t8, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:211:15  */
  assign n184_o = {1'b0, s7_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:211:23  */
  assign n185_o = {n184_o, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:211:31  */
  assign n186_o = ~d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:211:28  */
  assign n187_o = {n185_o, n186_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:211:39  */
  assign n189_o = {n187_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:212:21  */
  assign n190_o = t8s_h - u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:212:26  */
  assign n191_o = d8 ? n190_o : n192_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:213:20  */
  assign n192_o = t8s_h + u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:214:15  */
  assign n193_o = t10_h[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:215:16  */
  assign n194_o = {s7_d1, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:216:17  */
  assign n195_o = t9[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:216:11  */
  assign n196_o = ~n195_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:217:13  */
  assign n197_o = {s8, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:218:12  */
  assign n198_o = mr[8:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:219:15  */
  assign n199_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:220:39  */
  assign n201_o = {7'b0000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:220:16  */
  assign n202_o = fr + n201_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:221:19  */
  assign n203_o = {ern1_d2, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:224:21  */
  assign n206_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:225:21  */
  assign n209_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:226:21  */
  assign n212_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:227:21  */
  assign n215_o = xsx == 3'b001;
  assign n217_o = {n215_o, n212_o, n209_o, n206_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:223:4  */
  always @*
    case (n217_o)
      4'b1000: n218_o = 3'b001;
      4'b0100: n218_o = 3'b000;
      4'b0010: n218_o = 3'b100;
      4'b0001: n218_o = 3'b010;
      default: n218_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:229:16  */
  assign n219_o = {xsr_d2, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n220_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n221_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n222_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n223_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n224_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n225_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n226_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n227_q <= d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n228_q <= t7s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n229_q <= t7s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n230_q <= u7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n231_q <= s7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n232_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_8.vhdl:110:10  */
  always @(posedge clk)
    n233_q <= xsr_d1;
endmodule

