module fsqrt#(parameter ID=1)
  (input  clk,
   input  [33:0] X,
   output [33:0] R);
  wire [22:0] fracx;
  wire [7:0] ern0;
  wire [2:0] xsx;
  wire [7:0] ern1;
  wire [7:0] ern1_d1;
  wire [7:0] ern1_d2;
  wire [7:0] ern1_d3;
  wire [7:0] ern1_d4;
  wire [7:0] ern1_d5;
  wire [7:0] ern1_d6;
  wire [7:0] ern1_d7;
  wire [26:0] fracxnorm;
  wire [1:0] s0;
  wire [26:0] t1;
  wire d1;
  wire [27:0] t1s;
  wire [5:0] t1s_h;
  wire [21:0] t1s_l;
  wire [5:0] u1;
  wire [5:0] t3_h;
  wire [26:0] t2;
  wire [2:0] s1;
  wire d2;
  wire [27:0] t2s;
  wire [6:0] t2s_h;
  wire [20:0] t2s_l;
  wire [6:0] u2;
  wire [6:0] t4_h;
  wire [26:0] t3;
  wire [3:0] s2;
  wire d3;
  wire d3_d1;
  wire [27:0] t3s;
  wire [7:0] t3s_h;
  wire [7:0] t3s_h_d1;
  wire [19:0] t3s_l;
  wire [19:0] t3s_l_d1;
  wire [7:0] u3;
  wire [7:0] u3_d1;
  wire [7:0] t5_h;
  wire [26:0] t4;
  wire [4:0] s3;
  wire [4:0] s3_d1;
  wire d4;
  wire [27:0] t4s;
  wire [8:0] t4s_h;
  wire [18:0] t4s_l;
  wire [8:0] u4;
  wire [8:0] t6_h;
  wire [26:0] t5;
  wire [5:0] s4;
  wire d5;
  wire [27:0] t5s;
  wire [9:0] t5s_h;
  wire [17:0] t5s_l;
  wire [9:0] u5;
  wire [9:0] t7_h;
  wire [26:0] t6;
  wire [6:0] s5;
  wire d6;
  wire [27:0] t6s;
  wire [10:0] t6s_h;
  wire [16:0] t6s_l;
  wire [10:0] u6;
  wire [10:0] t8_h;
  wire [26:0] t7;
  wire [7:0] s6;
  wire d7;
  wire d7_d1;
  wire [27:0] t7s;
  wire [11:0] t7s_h;
  wire [11:0] t7s_h_d1;
  wire [15:0] t7s_l;
  wire [15:0] t7s_l_d1;
  wire [11:0] u7;
  wire [11:0] u7_d1;
  wire [11:0] t9_h;
  wire [26:0] t8;
  wire [8:0] s7;
  wire [8:0] s7_d1;
  wire d8;
  wire [27:0] t8s;
  wire [12:0] t8s_h;
  wire [14:0] t8s_l;
  wire [12:0] u8;
  wire [12:0] t10_h;
  wire [26:0] t9;
  wire [9:0] s8;
  wire d9;
  wire [27:0] t9s;
  wire [13:0] t9s_h;
  wire [13:0] t9s_l;
  wire [13:0] u9;
  wire [13:0] t11_h;
  wire [26:0] t10;
  wire [10:0] s9;
  wire d10;
  wire d10_d1;
  wire [27:0] t10s;
  wire [14:0] t10s_h;
  wire [14:0] t10s_h_d1;
  wire [12:0] t10s_l;
  wire [12:0] t10s_l_d1;
  wire [14:0] u10;
  wire [14:0] u10_d1;
  wire [14:0] t12_h;
  wire [26:0] t11;
  wire [11:0] s10;
  wire [11:0] s10_d1;
  wire d11;
  wire [27:0] t11s;
  wire [15:0] t11s_h;
  wire [11:0] t11s_l;
  wire [15:0] u11;
  wire [15:0] t13_h;
  wire [26:0] t12;
  wire [12:0] s11;
  wire d12;
  wire [27:0] t12s;
  wire [16:0] t12s_h;
  wire [10:0] t12s_l;
  wire [16:0] u12;
  wire [16:0] t14_h;
  wire [26:0] t13;
  wire [13:0] s12;
  wire d13;
  wire d13_d1;
  wire [27:0] t13s;
  wire [17:0] t13s_h;
  wire [17:0] t13s_h_d1;
  wire [9:0] t13s_l;
  wire [9:0] t13s_l_d1;
  wire [17:0] u13;
  wire [17:0] u13_d1;
  wire [17:0] t15_h;
  wire [26:0] t14;
  wire [14:0] s13;
  wire [14:0] s13_d1;
  wire d14;
  wire [27:0] t14s;
  wire [18:0] t14s_h;
  wire [8:0] t14s_l;
  wire [18:0] u14;
  wire [18:0] t16_h;
  wire [26:0] t15;
  wire [15:0] s14;
  wire d15;
  wire [27:0] t15s;
  wire [19:0] t15s_h;
  wire [7:0] t15s_l;
  wire [19:0] u15;
  wire [19:0] t17_h;
  wire [26:0] t16;
  wire [16:0] s15;
  wire d16;
  wire d16_d1;
  wire [27:0] t16s;
  wire [20:0] t16s_h;
  wire [20:0] t16s_h_d1;
  wire [6:0] t16s_l;
  wire [6:0] t16s_l_d1;
  wire [20:0] u16;
  wire [20:0] u16_d1;
  wire [20:0] t18_h;
  wire [26:0] t17;
  wire [17:0] s16;
  wire [17:0] s16_d1;
  wire d17;
  wire [27:0] t17s;
  wire [21:0] t17s_h;
  wire [5:0] t17s_l;
  wire [21:0] u17;
  wire [21:0] t19_h;
  wire [26:0] t18;
  wire [18:0] s17;
  wire d18;
  wire [27:0] t18s;
  wire [22:0] t18s_h;
  wire [4:0] t18s_l;
  wire [22:0] u18;
  wire [22:0] t20_h;
  wire [26:0] t19;
  wire [19:0] s18;
  wire d19;
  wire d19_d1;
  wire [27:0] t19s;
  wire [23:0] t19s_h;
  wire [23:0] t19s_h_d1;
  wire [3:0] t19s_l;
  wire [3:0] t19s_l_d1;
  wire [23:0] u19;
  wire [23:0] u19_d1;
  wire [23:0] t21_h;
  wire [26:0] t20;
  wire [20:0] s19;
  wire [20:0] s19_d1;
  wire d20;
  wire [27:0] t20s;
  wire [24:0] t20s_h;
  wire [2:0] t20s_l;
  wire [24:0] u20;
  wire [24:0] t22_h;
  wire [26:0] t21;
  wire [21:0] s20;
  wire d21;
  wire [27:0] t21s;
  wire [25:0] t21s_h;
  wire [1:0] t21s_l;
  wire [25:0] u21;
  wire [25:0] t23_h;
  wire [26:0] t22;
  wire [22:0] s21;
  wire d22;
  wire d22_d1;
  wire [27:0] t22s;
  wire [26:0] t22s_h;
  wire [26:0] t22s_h_d1;
  wire t22s_l;
  wire t22s_l_d1;
  wire [26:0] u22;
  wire [26:0] u22_d1;
  wire [26:0] t24_h;
  wire [26:0] t23;
  wire [23:0] s22;
  wire [23:0] s22_d1;
  wire d23;
  wire [27:0] t23s;
  wire [27:0] t23s_h;
  wire [27:0] u23;
  wire [27:0] t25_h;
  wire [26:0] t24;
  wire [24:0] s23;
  wire d25;
  wire [25:0] mr;
  wire [22:0] fr;
  wire round;
  wire [22:0] frrnd;
  wire [30:0] rn2;
  wire [2:0] xsr;
  wire [2:0] xsr_d1;
  wire [2:0] xsr_d2;
  wire [2:0] xsr_d3;
  wire [2:0] xsr_d4;
  wire [2:0] xsr_d5;
  wire [2:0] xsr_d6;
  wire [2:0] xsr_d7;
  wire [22:0] n54_o;
  wire [6:0] n55_o;
  wire [7:0] n57_o;
  wire [2:0] n58_o;
  wire [7:0] n60_o;
  wire n61_o;
  wire [7:0] n62_o;
  wire [7:0] n63_o;
  wire [23:0] n65_o;
  wire [26:0] n67_o;
  wire n68_o;
  wire n69_o;
  wire [26:0] n70_o;
  wire [24:0] n72_o;
  wire [26:0] n74_o;
  wire [3:0] n76_o;
  wire [3:0] n78_o;
  wire [22:0] n79_o;
  wire [26:0] n80_o;
  wire n81_o;
  wire n82_o;
  wire [27:0] n84_o;
  wire [5:0] n85_o;
  wire [21:0] n86_o;
  wire [2:0] n88_o;
  wire [3:0] n89_o;
  wire n90_o;
  wire [4:0] n91_o;
  wire [5:0] n93_o;
  wire [5:0] n94_o;
  wire [5:0] n95_o;
  wire [5:0] n96_o;
  wire [4:0] n97_o;
  wire [26:0] n98_o;
  wire [2:0] n99_o;
  wire n100_o;
  wire n101_o;
  wire [27:0] n103_o;
  wire [6:0] n104_o;
  wire [20:0] n105_o;
  wire [3:0] n107_o;
  wire [4:0] n108_o;
  wire n109_o;
  wire [5:0] n110_o;
  wire [6:0] n112_o;
  wire [6:0] n113_o;
  wire [6:0] n114_o;
  wire [6:0] n115_o;
  wire [5:0] n116_o;
  wire [26:0] n117_o;
  wire [3:0] n118_o;
  wire n119_o;
  wire n120_o;
  wire [27:0] n122_o;
  wire [7:0] n123_o;
  wire [19:0] n124_o;
  wire [4:0] n126_o;
  wire [5:0] n127_o;
  wire n128_o;
  wire [6:0] n129_o;
  wire [7:0] n131_o;
  wire [7:0] n132_o;
  wire [7:0] n133_o;
  wire [7:0] n134_o;
  wire [6:0] n135_o;
  wire [26:0] n136_o;
  wire [4:0] n137_o;
  wire n138_o;
  wire n139_o;
  wire [27:0] n141_o;
  wire [8:0] n142_o;
  wire [18:0] n143_o;
  wire [5:0] n145_o;
  wire [6:0] n146_o;
  wire n147_o;
  wire [7:0] n148_o;
  wire [8:0] n150_o;
  wire [8:0] n151_o;
  wire [8:0] n152_o;
  wire [8:0] n153_o;
  wire [7:0] n154_o;
  wire [26:0] n155_o;
  wire [5:0] n156_o;
  wire n157_o;
  wire n158_o;
  wire [27:0] n160_o;
  wire [9:0] n161_o;
  wire [17:0] n162_o;
  wire [6:0] n164_o;
  wire [7:0] n165_o;
  wire n166_o;
  wire [8:0] n167_o;
  wire [9:0] n169_o;
  wire [9:0] n170_o;
  wire [9:0] n171_o;
  wire [9:0] n172_o;
  wire [8:0] n173_o;
  wire [26:0] n174_o;
  wire [6:0] n175_o;
  wire n176_o;
  wire n177_o;
  wire [27:0] n179_o;
  wire [10:0] n180_o;
  wire [16:0] n181_o;
  wire [7:0] n183_o;
  wire [8:0] n184_o;
  wire n185_o;
  wire [9:0] n186_o;
  wire [10:0] n188_o;
  wire [10:0] n189_o;
  wire [10:0] n190_o;
  wire [10:0] n191_o;
  wire [9:0] n192_o;
  wire [26:0] n193_o;
  wire [7:0] n194_o;
  wire n195_o;
  wire n196_o;
  wire [27:0] n198_o;
  wire [11:0] n199_o;
  wire [15:0] n200_o;
  wire [8:0] n202_o;
  wire [9:0] n203_o;
  wire n204_o;
  wire [10:0] n205_o;
  wire [11:0] n207_o;
  wire [11:0] n208_o;
  wire [11:0] n209_o;
  wire [11:0] n210_o;
  wire [10:0] n211_o;
  wire [26:0] n212_o;
  wire [8:0] n213_o;
  wire n214_o;
  wire n215_o;
  wire [27:0] n217_o;
  wire [12:0] n218_o;
  wire [14:0] n219_o;
  wire [9:0] n221_o;
  wire [10:0] n222_o;
  wire n223_o;
  wire [11:0] n224_o;
  wire [12:0] n226_o;
  wire [12:0] n227_o;
  wire [12:0] n228_o;
  wire [12:0] n229_o;
  wire [11:0] n230_o;
  wire [26:0] n231_o;
  wire [9:0] n232_o;
  wire n233_o;
  wire n234_o;
  wire [27:0] n236_o;
  wire [13:0] n237_o;
  wire [13:0] n238_o;
  wire [10:0] n240_o;
  wire [11:0] n241_o;
  wire n242_o;
  wire [12:0] n243_o;
  wire [13:0] n245_o;
  wire [13:0] n246_o;
  wire [13:0] n247_o;
  wire [13:0] n248_o;
  wire [12:0] n249_o;
  wire [26:0] n250_o;
  wire [10:0] n251_o;
  wire n252_o;
  wire n253_o;
  wire [27:0] n255_o;
  wire [14:0] n256_o;
  wire [12:0] n257_o;
  wire [11:0] n259_o;
  wire [12:0] n260_o;
  wire n261_o;
  wire [13:0] n262_o;
  wire [14:0] n264_o;
  wire [14:0] n265_o;
  wire [14:0] n266_o;
  wire [14:0] n267_o;
  wire [13:0] n268_o;
  wire [26:0] n269_o;
  wire [11:0] n270_o;
  wire n271_o;
  wire n272_o;
  wire [27:0] n274_o;
  wire [15:0] n275_o;
  wire [11:0] n276_o;
  wire [12:0] n278_o;
  wire [13:0] n279_o;
  wire n280_o;
  wire [14:0] n281_o;
  wire [15:0] n283_o;
  wire [15:0] n284_o;
  wire [15:0] n285_o;
  wire [15:0] n286_o;
  wire [14:0] n287_o;
  wire [26:0] n288_o;
  wire [12:0] n289_o;
  wire n290_o;
  wire n291_o;
  wire [27:0] n293_o;
  wire [16:0] n294_o;
  wire [10:0] n295_o;
  wire [13:0] n297_o;
  wire [14:0] n298_o;
  wire n299_o;
  wire [15:0] n300_o;
  wire [16:0] n302_o;
  wire [16:0] n303_o;
  wire [16:0] n304_o;
  wire [16:0] n305_o;
  wire [15:0] n306_o;
  wire [26:0] n307_o;
  wire [13:0] n308_o;
  wire n309_o;
  wire n310_o;
  wire [27:0] n312_o;
  wire [17:0] n313_o;
  wire [9:0] n314_o;
  wire [14:0] n316_o;
  wire [15:0] n317_o;
  wire n318_o;
  wire [16:0] n319_o;
  wire [17:0] n321_o;
  wire [17:0] n322_o;
  wire [17:0] n323_o;
  wire [17:0] n324_o;
  wire [16:0] n325_o;
  wire [26:0] n326_o;
  wire [14:0] n327_o;
  wire n328_o;
  wire n329_o;
  wire [27:0] n331_o;
  wire [18:0] n332_o;
  wire [8:0] n333_o;
  wire [15:0] n335_o;
  wire [16:0] n336_o;
  wire n337_o;
  wire [17:0] n338_o;
  wire [18:0] n340_o;
  wire [18:0] n341_o;
  wire [18:0] n342_o;
  wire [18:0] n343_o;
  wire [17:0] n344_o;
  wire [26:0] n345_o;
  wire [15:0] n346_o;
  wire n347_o;
  wire n348_o;
  wire [27:0] n350_o;
  wire [19:0] n351_o;
  wire [7:0] n352_o;
  wire [16:0] n354_o;
  wire [17:0] n355_o;
  wire n356_o;
  wire [18:0] n357_o;
  wire [19:0] n359_o;
  wire [19:0] n360_o;
  wire [19:0] n361_o;
  wire [19:0] n362_o;
  wire [18:0] n363_o;
  wire [26:0] n364_o;
  wire [16:0] n365_o;
  wire n366_o;
  wire n367_o;
  wire [27:0] n369_o;
  wire [20:0] n370_o;
  wire [6:0] n371_o;
  wire [17:0] n373_o;
  wire [18:0] n374_o;
  wire n375_o;
  wire [19:0] n376_o;
  wire [20:0] n378_o;
  wire [20:0] n379_o;
  wire [20:0] n380_o;
  wire [20:0] n381_o;
  wire [19:0] n382_o;
  wire [26:0] n383_o;
  wire [17:0] n384_o;
  wire n385_o;
  wire n386_o;
  wire [27:0] n388_o;
  wire [21:0] n389_o;
  wire [5:0] n390_o;
  wire [18:0] n392_o;
  wire [19:0] n393_o;
  wire n394_o;
  wire [20:0] n395_o;
  wire [21:0] n397_o;
  wire [21:0] n398_o;
  wire [21:0] n399_o;
  wire [21:0] n400_o;
  wire [20:0] n401_o;
  wire [26:0] n402_o;
  wire [18:0] n403_o;
  wire n404_o;
  wire n405_o;
  wire [27:0] n407_o;
  wire [22:0] n408_o;
  wire [4:0] n409_o;
  wire [19:0] n411_o;
  wire [20:0] n412_o;
  wire n413_o;
  wire [21:0] n414_o;
  wire [22:0] n416_o;
  wire [22:0] n417_o;
  wire [22:0] n418_o;
  wire [22:0] n419_o;
  wire [21:0] n420_o;
  wire [26:0] n421_o;
  wire [19:0] n422_o;
  wire n423_o;
  wire n424_o;
  wire [27:0] n426_o;
  wire [23:0] n427_o;
  wire [3:0] n428_o;
  wire [20:0] n430_o;
  wire [21:0] n431_o;
  wire n432_o;
  wire [22:0] n433_o;
  wire [23:0] n435_o;
  wire [23:0] n436_o;
  wire [23:0] n437_o;
  wire [23:0] n438_o;
  wire [22:0] n439_o;
  wire [26:0] n440_o;
  wire [20:0] n441_o;
  wire n442_o;
  wire n443_o;
  wire [27:0] n445_o;
  wire [24:0] n446_o;
  wire [2:0] n447_o;
  wire [21:0] n449_o;
  wire [22:0] n450_o;
  wire n451_o;
  wire [23:0] n452_o;
  wire [24:0] n454_o;
  wire [24:0] n455_o;
  wire [24:0] n456_o;
  wire [24:0] n457_o;
  wire [23:0] n458_o;
  wire [26:0] n459_o;
  wire [21:0] n460_o;
  wire n461_o;
  wire n462_o;
  wire [27:0] n464_o;
  wire [25:0] n465_o;
  wire [1:0] n466_o;
  wire [22:0] n468_o;
  wire [23:0] n469_o;
  wire n470_o;
  wire [24:0] n471_o;
  wire [25:0] n473_o;
  wire [25:0] n474_o;
  wire [25:0] n475_o;
  wire [25:0] n476_o;
  wire [24:0] n477_o;
  wire [26:0] n478_o;
  wire [22:0] n479_o;
  wire n480_o;
  wire n481_o;
  wire [27:0] n483_o;
  wire [26:0] n484_o;
  wire n485_o;
  wire [23:0] n487_o;
  wire [24:0] n488_o;
  wire n489_o;
  wire [25:0] n490_o;
  wire [26:0] n492_o;
  wire [26:0] n493_o;
  wire [26:0] n494_o;
  wire [26:0] n495_o;
  wire [25:0] n496_o;
  wire [26:0] n497_o;
  wire [23:0] n498_o;
  wire n499_o;
  wire n500_o;
  wire [27:0] n502_o;
  wire [24:0] n504_o;
  wire [25:0] n505_o;
  wire n506_o;
  wire [26:0] n507_o;
  wire [27:0] n509_o;
  wire [27:0] n510_o;
  wire [27:0] n511_o;
  wire [27:0] n512_o;
  wire [26:0] n513_o;
  wire [24:0] n514_o;
  wire n515_o;
  wire n516_o;
  wire [25:0] n517_o;
  wire [22:0] n518_o;
  wire n519_o;
  wire [22:0] n521_o;
  wire [22:0] n522_o;
  wire [30:0] n523_o;
  wire n526_o;
  wire n529_o;
  wire n532_o;
  wire n535_o;
  wire [3:0] n537_o;
  reg [2:0] n538_o;
  wire [33:0] n539_o;
  reg [7:0] n540_q;
  reg [7:0] n541_q;
  reg [7:0] n542_q;
  reg [7:0] n543_q;
  reg [7:0] n544_q;
  reg [7:0] n545_q;
  reg [7:0] n546_q;
  reg n547_q;
  reg [7:0] n548_q;
  reg [19:0] n549_q;
  reg [7:0] n550_q;
  reg [4:0] n551_q;
  reg n552_q;
  reg [11:0] n553_q;
  reg [15:0] n554_q;
  reg [11:0] n555_q;
  reg [8:0] n556_q;
  reg n557_q;
  reg [14:0] n558_q;
  reg [12:0] n559_q;
  reg [14:0] n560_q;
  reg [11:0] n561_q;
  reg n562_q;
  reg [17:0] n563_q;
  reg [9:0] n564_q;
  reg [17:0] n565_q;
  reg [14:0] n566_q;
  reg n567_q;
  reg [20:0] n568_q;
  reg [6:0] n569_q;
  reg [20:0] n570_q;
  reg [17:0] n571_q;
  reg n572_q;
  reg [23:0] n573_q;
  reg [3:0] n574_q;
  reg [23:0] n575_q;
  reg [20:0] n576_q;
  reg n577_q;
  reg [26:0] n578_q;
  reg n579_q;
  reg [26:0] n580_q;
  reg [23:0] n581_q;
  reg [2:0] n582_q;
  reg [2:0] n583_q;
  reg [2:0] n584_q;
  reg [2:0] n585_q;
  reg [2:0] n586_q;
  reg [2:0] n587_q;
  reg [2:0] n588_q;
  assign R = n539_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:30:8  */
  assign fracx = n54_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:31:8  */
  assign ern0 = n57_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:32:8  */
  assign xsx = n58_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:8  */
  assign ern1 = n63_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:14  */
  assign ern1_d1 = n540_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:23  */
  assign ern1_d2 = n541_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:32  */
  assign ern1_d3 = n542_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:41  */
  assign ern1_d4 = n543_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:50  */
  assign ern1_d5 = n544_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:59  */
  assign ern1_d6 = n545_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:33:68  */
  assign ern1_d7 = n546_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:34:8  */
  assign fracxnorm = n70_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:35:8  */
  assign s0 = 2'b01; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:36:8  */
  assign t1 = n80_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:37:8  */
  assign d1 = n82_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:38:8  */
  assign t1s = n84_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:39:8  */
  assign t1s_h = n85_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:40:8  */
  assign t1s_l = n86_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:41:8  */
  assign u1 = n93_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:42:8  */
  assign t3_h = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:43:8  */
  assign t2 = n98_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:44:8  */
  assign s1 = n99_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:45:8  */
  assign d2 = n101_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:46:8  */
  assign t2s = n103_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:47:8  */
  assign t2s_h = n104_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:48:8  */
  assign t2s_l = n105_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:49:8  */
  assign u2 = n112_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:50:8  */
  assign t4_h = n114_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:51:8  */
  assign t3 = n117_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:52:8  */
  assign s2 = n118_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:53:8  */
  assign d3 = n120_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:53:12  */
  assign d3_d1 = n547_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:54:8  */
  assign t3s = n122_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:55:8  */
  assign t3s_h = n123_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:55:15  */
  assign t3s_h_d1 = n548_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:56:8  */
  assign t3s_l = n124_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:56:15  */
  assign t3s_l_d1 = n549_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:57:8  */
  assign u3 = n131_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:57:12  */
  assign u3_d1 = n550_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:58:8  */
  assign t5_h = n133_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:59:8  */
  assign t4 = n136_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:60:8  */
  assign s3 = n137_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:60:12  */
  assign s3_d1 = n551_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:61:8  */
  assign d4 = n139_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:62:8  */
  assign t4s = n141_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:63:8  */
  assign t4s_h = n142_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:64:8  */
  assign t4s_l = n143_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:65:8  */
  assign u4 = n150_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:66:8  */
  assign t6_h = n152_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:67:8  */
  assign t5 = n155_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:68:8  */
  assign s4 = n156_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:69:8  */
  assign d5 = n158_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:70:8  */
  assign t5s = n160_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:71:8  */
  assign t5s_h = n161_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:72:8  */
  assign t5s_l = n162_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:73:8  */
  assign u5 = n169_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:74:8  */
  assign t7_h = n171_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:75:8  */
  assign t6 = n174_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:76:8  */
  assign s5 = n175_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:77:8  */
  assign d6 = n177_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:78:8  */
  assign t6s = n179_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:79:8  */
  assign t6s_h = n180_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:80:8  */
  assign t6s_l = n181_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:81:8  */
  assign u6 = n188_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:82:8  */
  assign t8_h = n190_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:83:8  */
  assign t7 = n193_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:84:8  */
  assign s6 = n194_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:85:8  */
  assign d7 = n196_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:85:12  */
  assign d7_d1 = n552_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:86:8  */
  assign t7s = n198_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:87:8  */
  assign t7s_h = n199_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:87:15  */
  assign t7s_h_d1 = n553_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:88:8  */
  assign t7s_l = n200_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:88:15  */
  assign t7s_l_d1 = n554_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:89:8  */
  assign u7 = n207_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:89:12  */
  assign u7_d1 = n555_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:90:8  */
  assign t9_h = n209_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:91:8  */
  assign t8 = n212_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:92:8  */
  assign s7 = n213_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:92:12  */
  assign s7_d1 = n556_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:93:8  */
  assign d8 = n215_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:94:8  */
  assign t8s = n217_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:95:8  */
  assign t8s_h = n218_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:96:8  */
  assign t8s_l = n219_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:97:8  */
  assign u8 = n226_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:98:8  */
  assign t10_h = n228_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:99:8  */
  assign t9 = n231_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:100:8  */
  assign s8 = n232_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:101:8  */
  assign d9 = n234_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:102:8  */
  assign t9s = n236_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:103:8  */
  assign t9s_h = n237_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:104:8  */
  assign t9s_l = n238_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:105:8  */
  assign u9 = n245_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:106:8  */
  assign t11_h = n247_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:107:8  */
  assign t10 = n250_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:108:8  */
  assign s9 = n251_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:109:8  */
  assign d10 = n253_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:109:13  */
  assign d10_d1 = n557_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:110:8  */
  assign t10s = n255_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:111:8  */
  assign t10s_h = n256_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:111:16  */
  assign t10s_h_d1 = n558_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:112:8  */
  assign t10s_l = n257_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:112:16  */
  assign t10s_l_d1 = n559_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:113:8  */
  assign u10 = n264_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:113:13  */
  assign u10_d1 = n560_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:114:8  */
  assign t12_h = n266_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:115:8  */
  assign t11 = n269_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:116:8  */
  assign s10 = n270_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:116:13  */
  assign s10_d1 = n561_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:117:8  */
  assign d11 = n272_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:118:8  */
  assign t11s = n274_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:119:8  */
  assign t11s_h = n275_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:120:8  */
  assign t11s_l = n276_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:121:8  */
  assign u11 = n283_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:122:8  */
  assign t13_h = n285_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:123:8  */
  assign t12 = n288_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:124:8  */
  assign s11 = n289_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:125:8  */
  assign d12 = n291_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:126:8  */
  assign t12s = n293_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:127:8  */
  assign t12s_h = n294_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:128:8  */
  assign t12s_l = n295_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:129:8  */
  assign u12 = n302_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:130:8  */
  assign t14_h = n304_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:131:8  */
  assign t13 = n307_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:132:8  */
  assign s12 = n308_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:133:8  */
  assign d13 = n310_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:133:13  */
  assign d13_d1 = n562_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:134:8  */
  assign t13s = n312_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:135:8  */
  assign t13s_h = n313_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:135:16  */
  assign t13s_h_d1 = n563_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:136:8  */
  assign t13s_l = n314_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:136:16  */
  assign t13s_l_d1 = n564_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:137:8  */
  assign u13 = n321_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:137:13  */
  assign u13_d1 = n565_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:138:8  */
  assign t15_h = n323_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:139:8  */
  assign t14 = n326_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:140:8  */
  assign s13 = n327_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:140:13  */
  assign s13_d1 = n566_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:141:8  */
  assign d14 = n329_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:142:8  */
  assign t14s = n331_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:143:8  */
  assign t14s_h = n332_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:144:8  */
  assign t14s_l = n333_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:145:8  */
  assign u14 = n340_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:146:8  */
  assign t16_h = n342_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:147:8  */
  assign t15 = n345_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:148:8  */
  assign s14 = n346_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:149:8  */
  assign d15 = n348_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:150:8  */
  assign t15s = n350_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:151:8  */
  assign t15s_h = n351_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:152:8  */
  assign t15s_l = n352_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:153:8  */
  assign u15 = n359_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:154:8  */
  assign t17_h = n361_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:155:8  */
  assign t16 = n364_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:156:8  */
  assign s15 = n365_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:157:8  */
  assign d16 = n367_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:157:13  */
  assign d16_d1 = n567_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:158:8  */
  assign t16s = n369_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:159:8  */
  assign t16s_h = n370_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:159:16  */
  assign t16s_h_d1 = n568_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:160:8  */
  assign t16s_l = n371_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:160:16  */
  assign t16s_l_d1 = n569_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:161:8  */
  assign u16 = n378_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:161:13  */
  assign u16_d1 = n570_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:162:8  */
  assign t18_h = n380_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:163:8  */
  assign t17 = n383_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:164:8  */
  assign s16 = n384_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:164:13  */
  assign s16_d1 = n571_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:165:8  */
  assign d17 = n386_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:166:8  */
  assign t17s = n388_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:167:8  */
  assign t17s_h = n389_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:168:8  */
  assign t17s_l = n390_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:169:8  */
  assign u17 = n397_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:170:8  */
  assign t19_h = n399_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:171:8  */
  assign t18 = n402_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:172:8  */
  assign s17 = n403_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:173:8  */
  assign d18 = n405_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:174:8  */
  assign t18s = n407_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:175:8  */
  assign t18s_h = n408_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:176:8  */
  assign t18s_l = n409_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:177:8  */
  assign u18 = n416_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:178:8  */
  assign t20_h = n418_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:179:8  */
  assign t19 = n421_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:180:8  */
  assign s18 = n422_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:181:8  */
  assign d19 = n424_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:181:13  */
  assign d19_d1 = n572_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:182:8  */
  assign t19s = n426_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:183:8  */
  assign t19s_h = n427_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:183:16  */
  assign t19s_h_d1 = n573_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:184:8  */
  assign t19s_l = n428_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:184:16  */
  assign t19s_l_d1 = n574_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:185:8  */
  assign u19 = n435_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:185:13  */
  assign u19_d1 = n575_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:186:8  */
  assign t21_h = n437_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:187:8  */
  assign t20 = n440_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:188:8  */
  assign s19 = n441_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:188:13  */
  assign s19_d1 = n576_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:189:8  */
  assign d20 = n443_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:190:8  */
  assign t20s = n445_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:191:8  */
  assign t20s_h = n446_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:192:8  */
  assign t20s_l = n447_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:193:8  */
  assign u20 = n454_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:194:8  */
  assign t22_h = n456_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:195:8  */
  assign t21 = n459_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:196:8  */
  assign s20 = n460_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:197:8  */
  assign d21 = n462_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:198:8  */
  assign t21s = n464_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:199:8  */
  assign t21s_h = n465_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:200:8  */
  assign t21s_l = n466_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:201:8  */
  assign u21 = n473_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:202:8  */
  assign t23_h = n475_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:203:8  */
  assign t22 = n478_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:204:8  */
  assign s21 = n479_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:205:8  */
  assign d22 = n481_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:205:13  */
  assign d22_d1 = n577_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:206:8  */
  assign t22s = n483_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:207:8  */
  assign t22s_h = n484_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:207:16  */
  assign t22s_h_d1 = n578_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:208:8  */
  assign t22s_l = n485_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:208:16  */
  assign t22s_l_d1 = n579_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:209:8  */
  assign u22 = n492_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:209:13  */
  assign u22_d1 = n580_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:210:8  */
  assign t24_h = n494_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:211:8  */
  assign t23 = n497_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:212:8  */
  assign s22 = n498_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:212:13  */
  assign s22_d1 = n581_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:213:8  */
  assign d23 = n500_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:515:18  */
  assign t23s = n502_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:215:8  */
  assign t23s_h = t23s; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:216:8  */
  assign u23 = n509_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:217:8  */
  assign t25_h = n511_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:218:8  */
  assign t24 = n513_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:219:8  */
  assign s23 = n514_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:220:8  */
  assign d25 = n516_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:221:8  */
  assign mr = n517_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:222:8  */
  assign fr = n518_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:223:8  */
  assign round = n519_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:224:8  */
  assign frrnd = n522_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:225:8  */
  assign rn2 = n523_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:8  */
  assign xsr = n538_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:13  */
  assign xsr_d1 = n582_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:21  */
  assign xsr_d2 = n583_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:29  */
  assign xsr_d3 = n584_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:37  */
  assign xsr_d4 = n585_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:45  */
  assign xsr_d5 = n586_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:53  */
  assign xsr_d6 = n587_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:226:61  */
  assign xsr_d7 = n588_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:282:14  */
  assign n54_o = X[22:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:283:19  */
  assign n55_o = X[30:24];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:283:16  */
  assign n57_o = {1'b0, n55_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:284:12  */
  assign n58_o = X[33:31];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:285:17  */
  assign n60_o = ern0 + 8'b00111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:285:51  */
  assign n61_o = X[23];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:285:48  */
  assign n62_o = {7'b0, n61_o};  //  uext
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:285:48  */
  assign n63_o = n60_o + n62_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:286:21  */
  assign n65_o = {1'b1, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:286:29  */
  assign n67_o = {n65_o, 3'b000};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:286:43  */
  assign n68_o = X[23];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:286:48  */
  assign n69_o = ~n68_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:286:37  */
  assign n70_o = n69_o ? n67_o : n74_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:287:15  */
  assign n72_o = {2'b01, fracx};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:287:22  */
  assign n74_o = {n72_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:289:29  */
  assign n76_o = fracxnorm[26:23];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:289:18  */
  assign n78_o = 4'b0111 + n76_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:289:56  */
  assign n79_o = fracxnorm[22:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:289:45  */
  assign n80_o = {n78_o, n79_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:293:16  */
  assign n81_o = t1[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:293:10  */
  assign n82_o = ~n81_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:294:14  */
  assign n84_o = {t1, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:295:16  */
  assign n85_o = t1s[27:22];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:296:16  */
  assign n86_o = t1s[21:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:297:15  */
  assign n88_o = {1'b0, s0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:297:20  */
  assign n89_o = {n88_o, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:297:28  */
  assign n90_o = ~d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:297:25  */
  assign n91_o = {n89_o, n90_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:297:36  */
  assign n93_o = {n91_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:298:20  */
  assign n94_o = t1s_h - u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:298:25  */
  assign n95_o = d1 ? n94_o : n96_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:299:20  */
  assign n96_o = t1s_h + u1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:300:14  */
  assign n97_o = t3_h[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:300:27  */
  assign n98_o = {n97_o, t1s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:301:13  */
  assign n99_o = {s0, d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:303:16  */
  assign n100_o = t2[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:303:10  */
  assign n101_o = ~n100_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:304:14  */
  assign n103_o = {t2, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:305:16  */
  assign n104_o = t2s[27:21];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:306:16  */
  assign n105_o = t2s[20:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:307:15  */
  assign n107_o = {1'b0, s1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:307:20  */
  assign n108_o = {n107_o, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:307:28  */
  assign n109_o = ~d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:307:25  */
  assign n110_o = {n108_o, n109_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:307:36  */
  assign n112_o = {n110_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:308:20  */
  assign n113_o = t2s_h - u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:308:25  */
  assign n114_o = d2 ? n113_o : n115_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:309:20  */
  assign n115_o = t2s_h + u2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:310:14  */
  assign n116_o = t4_h[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:310:27  */
  assign n117_o = {n116_o, t2s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:311:13  */
  assign n118_o = {s1, d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:313:16  */
  assign n119_o = t3[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:313:10  */
  assign n120_o = ~n119_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:314:14  */
  assign n122_o = {t3, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:315:16  */
  assign n123_o = t3s[27:20];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:316:16  */
  assign n124_o = t3s[19:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:317:15  */
  assign n126_o = {1'b0, s2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:317:20  */
  assign n127_o = {n126_o, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:317:28  */
  assign n128_o = ~d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:317:25  */
  assign n129_o = {n127_o, n128_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:317:36  */
  assign n131_o = {n129_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:318:23  */
  assign n132_o = t3s_h_d1 - u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:318:31  */
  assign n133_o = d3_d1 ? n132_o : n134_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:319:23  */
  assign n134_o = t3s_h_d1 + u3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:320:14  */
  assign n135_o = t5_h[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:320:27  */
  assign n136_o = {n135_o, t3s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:321:13  */
  assign n137_o = {s2, d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:323:16  */
  assign n138_o = t4[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:323:10  */
  assign n139_o = ~n138_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:324:14  */
  assign n141_o = {t4, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:325:16  */
  assign n142_o = t4s[27:19];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:326:16  */
  assign n143_o = t4s[18:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:327:15  */
  assign n145_o = {1'b0, s3_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:327:23  */
  assign n146_o = {n145_o, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:327:31  */
  assign n147_o = ~d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:327:28  */
  assign n148_o = {n146_o, n147_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:327:39  */
  assign n150_o = {n148_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:328:20  */
  assign n151_o = t4s_h - u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:328:25  */
  assign n152_o = d4 ? n151_o : n153_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:329:20  */
  assign n153_o = t4s_h + u4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:330:14  */
  assign n154_o = t6_h[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:330:27  */
  assign n155_o = {n154_o, t4s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:331:16  */
  assign n156_o = {s3_d1, d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:333:16  */
  assign n157_o = t5[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:333:10  */
  assign n158_o = ~n157_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:334:14  */
  assign n160_o = {t5, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:335:16  */
  assign n161_o = t5s[27:18];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:336:16  */
  assign n162_o = t5s[17:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:337:15  */
  assign n164_o = {1'b0, s4};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:337:20  */
  assign n165_o = {n164_o, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:337:28  */
  assign n166_o = ~d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:337:25  */
  assign n167_o = {n165_o, n166_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:337:36  */
  assign n169_o = {n167_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:338:20  */
  assign n170_o = t5s_h - u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:338:25  */
  assign n171_o = d5 ? n170_o : n172_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:339:20  */
  assign n172_o = t5s_h + u5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:340:14  */
  assign n173_o = t7_h[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:340:27  */
  assign n174_o = {n173_o, t5s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:341:13  */
  assign n175_o = {s4, d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:343:16  */
  assign n176_o = t6[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:343:10  */
  assign n177_o = ~n176_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:344:14  */
  assign n179_o = {t6, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:345:16  */
  assign n180_o = t6s[27:17];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:346:16  */
  assign n181_o = t6s[16:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:347:15  */
  assign n183_o = {1'b0, s5};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:347:20  */
  assign n184_o = {n183_o, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:347:28  */
  assign n185_o = ~d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:347:25  */
  assign n186_o = {n184_o, n185_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:347:36  */
  assign n188_o = {n186_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:348:20  */
  assign n189_o = t6s_h - u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:348:25  */
  assign n190_o = d6 ? n189_o : n191_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:349:20  */
  assign n191_o = t6s_h + u6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:350:14  */
  assign n192_o = t8_h[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:350:27  */
  assign n193_o = {n192_o, t6s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:351:13  */
  assign n194_o = {s5, d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:353:16  */
  assign n195_o = t7[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:353:10  */
  assign n196_o = ~n195_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:354:14  */
  assign n198_o = {t7, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:355:16  */
  assign n199_o = t7s[27:16];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:356:16  */
  assign n200_o = t7s[15:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:357:15  */
  assign n202_o = {1'b0, s6};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:357:20  */
  assign n203_o = {n202_o, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:357:28  */
  assign n204_o = ~d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:357:25  */
  assign n205_o = {n203_o, n204_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:357:36  */
  assign n207_o = {n205_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:358:23  */
  assign n208_o = t7s_h_d1 - u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:358:31  */
  assign n209_o = d7_d1 ? n208_o : n210_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:359:23  */
  assign n210_o = t7s_h_d1 + u7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:360:14  */
  assign n211_o = t9_h[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:360:28  */
  assign n212_o = {n211_o, t7s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:361:13  */
  assign n213_o = {s6, d7};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:363:16  */
  assign n214_o = t8[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:363:10  */
  assign n215_o = ~n214_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:364:14  */
  assign n217_o = {t8, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:365:16  */
  assign n218_o = t8s[27:15];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:366:16  */
  assign n219_o = t8s[14:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:367:15  */
  assign n221_o = {1'b0, s7_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:367:23  */
  assign n222_o = {n221_o, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:367:31  */
  assign n223_o = ~d8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:367:28  */
  assign n224_o = {n222_o, n223_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:367:39  */
  assign n226_o = {n224_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:368:21  */
  assign n227_o = t8s_h - u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:368:26  */
  assign n228_o = d8 ? n227_o : n229_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:369:20  */
  assign n229_o = t8s_h + u8;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:370:15  */
  assign n230_o = t10_h[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:370:29  */
  assign n231_o = {n230_o, t8s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:371:16  */
  assign n232_o = {s7_d1, d8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:373:16  */
  assign n233_o = t9[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:373:10  */
  assign n234_o = ~n233_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:374:14  */
  assign n236_o = {t9, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:375:16  */
  assign n237_o = t9s[27:14];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:376:16  */
  assign n238_o = t9s[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:377:15  */
  assign n240_o = {1'b0, s8};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:377:20  */
  assign n241_o = {n240_o, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:377:28  */
  assign n242_o = ~d9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:377:25  */
  assign n243_o = {n241_o, n242_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:377:36  */
  assign n245_o = {n243_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:378:21  */
  assign n246_o = t9s_h - u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:378:26  */
  assign n247_o = d9 ? n246_o : n248_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:379:20  */
  assign n248_o = t9s_h + u9;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:380:16  */
  assign n249_o = t11_h[12:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:380:30  */
  assign n250_o = {n249_o, t9s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:381:13  */
  assign n251_o = {s8, d9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:383:18  */
  assign n252_o = t10[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:383:11  */
  assign n253_o = ~n252_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:384:16  */
  assign n255_o = {t10, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:385:18  */
  assign n256_o = t10s[27:13];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:386:18  */
  assign n257_o = t10s[12:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:387:16  */
  assign n259_o = {1'b0, s9};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:387:21  */
  assign n260_o = {n259_o, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:387:30  */
  assign n261_o = ~d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:387:27  */
  assign n262_o = {n260_o, n261_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:387:39  */
  assign n264_o = {n262_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:388:25  */
  assign n265_o = t10s_h_d1 - u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:388:34  */
  assign n266_o = d10_d1 ? n265_o : n267_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:389:24  */
  assign n267_o = t10s_h_d1 + u10_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:390:16  */
  assign n268_o = t12_h[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:390:30  */
  assign n269_o = {n268_o, t10s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:391:14  */
  assign n270_o = {s9, d10};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:393:18  */
  assign n271_o = t11[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:393:11  */
  assign n272_o = ~n271_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:394:16  */
  assign n274_o = {t11, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:395:18  */
  assign n275_o = t11s[27:12];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:396:18  */
  assign n276_o = t11s[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:397:16  */
  assign n278_o = {1'b0, s10_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:397:25  */
  assign n279_o = {n278_o, d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:397:34  */
  assign n280_o = ~d11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:397:31  */
  assign n281_o = {n279_o, n280_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:397:43  */
  assign n283_o = {n281_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:398:22  */
  assign n284_o = t11s_h - u11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:398:28  */
  assign n285_o = d11 ? n284_o : n286_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:399:21  */
  assign n286_o = t11s_h + u11;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:400:16  */
  assign n287_o = t13_h[14:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:400:30  */
  assign n288_o = {n287_o, t11s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:401:18  */
  assign n289_o = {s10_d1, d11};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:403:18  */
  assign n290_o = t12[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:403:11  */
  assign n291_o = ~n290_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:404:16  */
  assign n293_o = {t12, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:405:18  */
  assign n294_o = t12s[27:11];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:406:18  */
  assign n295_o = t12s[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:407:16  */
  assign n297_o = {1'b0, s11};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:407:22  */
  assign n298_o = {n297_o, d12};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:407:31  */
  assign n299_o = ~d12;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:407:28  */
  assign n300_o = {n298_o, n299_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:407:40  */
  assign n302_o = {n300_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:408:22  */
  assign n303_o = t12s_h - u12;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:408:28  */
  assign n304_o = d12 ? n303_o : n305_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:409:21  */
  assign n305_o = t12s_h + u12;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:410:16  */
  assign n306_o = t14_h[15:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:410:30  */
  assign n307_o = {n306_o, t12s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:411:15  */
  assign n308_o = {s11, d12};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:413:18  */
  assign n309_o = t13[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:413:11  */
  assign n310_o = ~n309_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:414:16  */
  assign n312_o = {t13, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:415:18  */
  assign n313_o = t13s[27:10];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:416:18  */
  assign n314_o = t13s[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:417:16  */
  assign n316_o = {1'b0, s12};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:417:22  */
  assign n317_o = {n316_o, d13};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:417:31  */
  assign n318_o = ~d13;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:417:28  */
  assign n319_o = {n317_o, n318_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:417:40  */
  assign n321_o = {n319_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:418:25  */
  assign n322_o = t13s_h_d1 - u13_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:418:34  */
  assign n323_o = d13_d1 ? n322_o : n324_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:419:24  */
  assign n324_o = t13s_h_d1 + u13_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:420:16  */
  assign n325_o = t15_h[16:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:420:30  */
  assign n326_o = {n325_o, t13s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:421:15  */
  assign n327_o = {s12, d13};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:423:18  */
  assign n328_o = t14[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:423:11  */
  assign n329_o = ~n328_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:424:16  */
  assign n331_o = {t14, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:425:18  */
  assign n332_o = t14s[27:9];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:426:18  */
  assign n333_o = t14s[8:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:427:16  */
  assign n335_o = {1'b0, s13_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:427:25  */
  assign n336_o = {n335_o, d14};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:427:34  */
  assign n337_o = ~d14;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:427:31  */
  assign n338_o = {n336_o, n337_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:427:43  */
  assign n340_o = {n338_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:428:22  */
  assign n341_o = t14s_h - u14;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:428:28  */
  assign n342_o = d14 ? n341_o : n343_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:429:21  */
  assign n343_o = t14s_h + u14;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:430:16  */
  assign n344_o = t16_h[17:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:430:30  */
  assign n345_o = {n344_o, t14s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:431:18  */
  assign n346_o = {s13_d1, d14};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:433:18  */
  assign n347_o = t15[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:433:11  */
  assign n348_o = ~n347_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:434:16  */
  assign n350_o = {t15, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:435:18  */
  assign n351_o = t15s[27:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:436:18  */
  assign n352_o = t15s[7:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:437:16  */
  assign n354_o = {1'b0, s14};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:437:22  */
  assign n355_o = {n354_o, d15};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:437:31  */
  assign n356_o = ~d15;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:437:28  */
  assign n357_o = {n355_o, n356_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:437:40  */
  assign n359_o = {n357_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:438:22  */
  assign n360_o = t15s_h - u15;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:438:28  */
  assign n361_o = d15 ? n360_o : n362_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:439:21  */
  assign n362_o = t15s_h + u15;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:440:16  */
  assign n363_o = t17_h[18:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:440:30  */
  assign n364_o = {n363_o, t15s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:441:15  */
  assign n365_o = {s14, d15};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:443:18  */
  assign n366_o = t16[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:443:11  */
  assign n367_o = ~n366_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:444:16  */
  assign n369_o = {t16, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:445:18  */
  assign n370_o = t16s[27:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:446:18  */
  assign n371_o = t16s[6:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:447:16  */
  assign n373_o = {1'b0, s15};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:447:22  */
  assign n374_o = {n373_o, d16};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:447:31  */
  assign n375_o = ~d16;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:447:28  */
  assign n376_o = {n374_o, n375_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:447:40  */
  assign n378_o = {n376_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:448:25  */
  assign n379_o = t16s_h_d1 - u16_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:448:34  */
  assign n380_o = d16_d1 ? n379_o : n381_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:449:24  */
  assign n381_o = t16s_h_d1 + u16_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:450:16  */
  assign n382_o = t18_h[19:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:450:30  */
  assign n383_o = {n382_o, t16s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:451:15  */
  assign n384_o = {s15, d16};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:453:18  */
  assign n385_o = t17[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:453:11  */
  assign n386_o = ~n385_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:454:16  */
  assign n388_o = {t17, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:455:18  */
  assign n389_o = t17s[27:6];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:456:18  */
  assign n390_o = t17s[5:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:457:16  */
  assign n392_o = {1'b0, s16_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:457:25  */
  assign n393_o = {n392_o, d17};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:457:34  */
  assign n394_o = ~d17;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:457:31  */
  assign n395_o = {n393_o, n394_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:457:43  */
  assign n397_o = {n395_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:458:22  */
  assign n398_o = t17s_h - u17;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:458:28  */
  assign n399_o = d17 ? n398_o : n400_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:459:21  */
  assign n400_o = t17s_h + u17;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:460:16  */
  assign n401_o = t19_h[20:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:460:30  */
  assign n402_o = {n401_o, t17s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:461:18  */
  assign n403_o = {s16_d1, d17};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:463:18  */
  assign n404_o = t18[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:463:11  */
  assign n405_o = ~n404_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:464:16  */
  assign n407_o = {t18, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:465:18  */
  assign n408_o = t18s[27:5];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:466:18  */
  assign n409_o = t18s[4:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:467:16  */
  assign n411_o = {1'b0, s17};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:467:22  */
  assign n412_o = {n411_o, d18};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:467:31  */
  assign n413_o = ~d18;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:467:28  */
  assign n414_o = {n412_o, n413_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:467:40  */
  assign n416_o = {n414_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:468:22  */
  assign n417_o = t18s_h - u18;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:468:28  */
  assign n418_o = d18 ? n417_o : n419_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:469:21  */
  assign n419_o = t18s_h + u18;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:470:16  */
  assign n420_o = t20_h[21:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:470:30  */
  assign n421_o = {n420_o, t18s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:471:15  */
  assign n422_o = {s17, d18};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:473:18  */
  assign n423_o = t19[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:473:11  */
  assign n424_o = ~n423_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:474:16  */
  assign n426_o = {t19, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:475:18  */
  assign n427_o = t19s[27:4];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:476:18  */
  assign n428_o = t19s[3:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:477:16  */
  assign n430_o = {1'b0, s18};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:477:22  */
  assign n431_o = {n430_o, d19};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:477:31  */
  assign n432_o = ~d19;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:477:28  */
  assign n433_o = {n431_o, n432_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:477:40  */
  assign n435_o = {n433_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:478:25  */
  assign n436_o = t19s_h_d1 - u19_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:478:34  */
  assign n437_o = d19_d1 ? n436_o : n438_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:479:24  */
  assign n438_o = t19s_h_d1 + u19_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:480:16  */
  assign n439_o = t21_h[22:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:480:30  */
  assign n440_o = {n439_o, t19s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:481:15  */
  assign n441_o = {s18, d19};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:483:18  */
  assign n442_o = t20[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:483:11  */
  assign n443_o = ~n442_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:484:16  */
  assign n445_o = {t20, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:485:18  */
  assign n446_o = t20s[27:3];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:486:18  */
  assign n447_o = t20s[2:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:487:16  */
  assign n449_o = {1'b0, s19_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:487:25  */
  assign n450_o = {n449_o, d20};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:487:34  */
  assign n451_o = ~d20;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:487:31  */
  assign n452_o = {n450_o, n451_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:487:43  */
  assign n454_o = {n452_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:488:22  */
  assign n455_o = t20s_h - u20;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:488:28  */
  assign n456_o = d20 ? n455_o : n457_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:489:21  */
  assign n457_o = t20s_h + u20;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:490:16  */
  assign n458_o = t22_h[23:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:490:30  */
  assign n459_o = {n458_o, t20s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:491:18  */
  assign n460_o = {s19_d1, d20};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:493:18  */
  assign n461_o = t21[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:493:11  */
  assign n462_o = ~n461_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:494:16  */
  assign n464_o = {t21, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:495:18  */
  assign n465_o = t21s[27:2];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:496:18  */
  assign n466_o = t21s[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:497:16  */
  assign n468_o = {1'b0, s20};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:497:22  */
  assign n469_o = {n468_o, d21};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:497:31  */
  assign n470_o = ~d21;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:497:28  */
  assign n471_o = {n469_o, n470_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:497:40  */
  assign n473_o = {n471_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:498:22  */
  assign n474_o = t21s_h - u21;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:498:28  */
  assign n475_o = d21 ? n474_o : n476_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:499:21  */
  assign n476_o = t21s_h + u21;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:500:16  */
  assign n477_o = t23_h[24:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:500:30  */
  assign n478_o = {n477_o, t21s_l};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:501:15  */
  assign n479_o = {s20, d21};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:503:18  */
  assign n480_o = t22[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:503:11  */
  assign n481_o = ~n480_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:504:16  */
  assign n483_o = {t22, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:505:18  */
  assign n484_o = t22s[27:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:506:18  */
  assign n485_o = t22s[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:507:16  */
  assign n487_o = {1'b0, s21};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:507:22  */
  assign n488_o = {n487_o, d22};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:507:31  */
  assign n489_o = ~d22;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:507:28  */
  assign n490_o = {n488_o, n489_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:507:40  */
  assign n492_o = {n490_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:508:25  */
  assign n493_o = t22s_h_d1 - u22_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:508:34  */
  assign n494_o = d22_d1 ? n493_o : n495_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:509:24  */
  assign n495_o = t22s_h_d1 + u22_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:510:16  */
  assign n496_o = t24_h[25:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:510:30  */
  assign n497_o = {n496_o, t22s_l_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:511:15  */
  assign n498_o = {s21, d22};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:513:18  */
  assign n499_o = t23[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:513:11  */
  assign n500_o = ~n499_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:514:16  */
  assign n502_o = {t23, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:516:16  */
  assign n504_o = {1'b0, s22_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:516:25  */
  assign n505_o = {n504_o, d23};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:516:34  */
  assign n506_o = ~d23;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:516:31  */
  assign n507_o = {n505_o, n506_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:516:43  */
  assign n509_o = {n507_o, 1'b1};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:517:22  */
  assign n510_o = t23s_h - u23;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:517:28  */
  assign n511_o = d23 ? n510_o : n512_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:518:21  */
  assign n512_o = t23s_h + u23;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:519:16  */
  assign n513_o = t25_h[26:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:520:18  */
  assign n514_o = {s22_d1, d23};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:521:18  */
  assign n515_o = t24[26];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:521:11  */
  assign n516_o = ~n515_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:522:14  */
  assign n517_o = {s23, d25};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:523:12  */
  assign n518_o = mr[23:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:524:15  */
  assign n519_o = mr[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:525:40  */
  assign n521_o = {22'b0000000000000000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:525:16  */
  assign n522_o = fr + n521_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:526:19  */
  assign n523_o = {ern1_d7, frrnd};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:529:21  */
  assign n526_o = xsx == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:530:21  */
  assign n529_o = xsx == 3'b100;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:531:21  */
  assign n532_o = xsx == 3'b000;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:532:21  */
  assign n535_o = xsx == 3'b001;
  assign n537_o = {n535_o, n532_o, n529_o, n526_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:528:4  */
  always @*
    case (n537_o)
      4'b1000: n538_o = 3'b001;
      4'b0100: n538_o = 3'b000;
      4'b0010: n538_o = 3'b100;
      4'b0001: n538_o = 3'b010;
      default: n538_o = 3'b110;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:534:16  */
  assign n539_o = {xsr_d7, rn2};
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n540_q <= ern1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n541_q <= ern1_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n542_q <= ern1_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n543_q <= ern1_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n544_q <= ern1_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n545_q <= ern1_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n546_q <= ern1_d6;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n547_q <= d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n548_q <= t3s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n549_q <= t3s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n550_q <= u3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n551_q <= s3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n552_q <= d7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n553_q <= t7s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n554_q <= t7s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n555_q <= u7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n556_q <= s7;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n557_q <= d10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n558_q <= t10s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n559_q <= t10s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n560_q <= u10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n561_q <= s10;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n562_q <= d13;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n563_q <= t13s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n564_q <= t13s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n565_q <= u13;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n566_q <= s13;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n567_q <= d16;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n568_q <= t16s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n569_q <= t16s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n570_q <= u16;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n571_q <= s16;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n572_q <= d19;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n573_q <= t19s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n574_q <= t19s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n575_q <= u19;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n576_q <= s19;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n577_q <= d22;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n578_q <= t22s_h;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n579_q <= t22s_l;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n580_q <= u22;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n581_q <= s22;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n582_q <= xsr;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n583_q <= xsr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n584_q <= xsr_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n585_q <= xsr_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n586_q <= xsr_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n587_q <= xsr_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/flopoco_fsqrt_8_23.vhdl:230:10  */
  always @(posedge clk)
    n588_q <= xsr_d6;
endmodule

