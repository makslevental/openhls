module selfunction_f300_uid4
  (input wire [8:0] x,
   output wire [2:0] y);
  wire [2:0] y0;
  wire [2:0] y1;
  wire n509_o;
  wire n512_o;
  wire n515_o;
  wire n518_o;
  wire n521_o;
  wire n524_o;
  wire n527_o;
  wire n530_o;
  wire n533_o;
  wire n536_o;
  wire n539_o;
  wire n542_o;
  wire n545_o;
  wire n548_o;
  wire n551_o;
  wire n554_o;
  wire n557_o;
  wire n560_o;
  wire n563_o;
  wire n566_o;
  wire n569_o;
  wire n572_o;
  wire n575_o;
  wire n578_o;
  wire n581_o;
  wire n584_o;
  wire n587_o;
  wire n590_o;
  wire n593_o;
  wire n596_o;
  wire n599_o;
  wire n602_o;
  wire n605_o;
  wire n608_o;
  wire n611_o;
  wire n614_o;
  wire n617_o;
  wire n620_o;
  wire n623_o;
  wire n626_o;
  wire n629_o;
  wire n632_o;
  wire n635_o;
  wire n638_o;
  wire n641_o;
  wire n644_o;
  wire n647_o;
  wire n650_o;
  wire n653_o;
  wire n656_o;
  wire n659_o;
  wire n662_o;
  wire n665_o;
  wire n668_o;
  wire n671_o;
  wire n674_o;
  wire n677_o;
  wire n680_o;
  wire n683_o;
  wire n686_o;
  wire n689_o;
  wire n692_o;
  wire n695_o;
  wire n698_o;
  wire n701_o;
  wire n704_o;
  wire n707_o;
  wire n710_o;
  wire n713_o;
  wire n716_o;
  wire n719_o;
  wire n722_o;
  wire n725_o;
  wire n728_o;
  wire n731_o;
  wire n734_o;
  wire n737_o;
  wire n740_o;
  wire n743_o;
  wire n746_o;
  wire n749_o;
  wire n752_o;
  wire n755_o;
  wire n758_o;
  wire n761_o;
  wire n764_o;
  wire n767_o;
  wire n770_o;
  wire n773_o;
  wire n776_o;
  wire n779_o;
  wire n782_o;
  wire n785_o;
  wire n788_o;
  wire n791_o;
  wire n794_o;
  wire n797_o;
  wire n800_o;
  wire n803_o;
  wire n806_o;
  wire n809_o;
  wire n812_o;
  wire n815_o;
  wire n818_o;
  wire n821_o;
  wire n824_o;
  wire n827_o;
  wire n830_o;
  wire n833_o;
  wire n836_o;
  wire n839_o;
  wire n842_o;
  wire n845_o;
  wire n848_o;
  wire n851_o;
  wire n854_o;
  wire n857_o;
  wire n860_o;
  wire n863_o;
  wire n866_o;
  wire n869_o;
  wire n872_o;
  wire n875_o;
  wire n878_o;
  wire n881_o;
  wire n884_o;
  wire n887_o;
  wire n890_o;
  wire n893_o;
  wire n896_o;
  wire n899_o;
  wire n902_o;
  wire n905_o;
  wire n908_o;
  wire n911_o;
  wire n914_o;
  wire n917_o;
  wire n920_o;
  wire n923_o;
  wire n926_o;
  wire n929_o;
  wire n932_o;
  wire n935_o;
  wire n938_o;
  wire n941_o;
  wire n944_o;
  wire n947_o;
  wire n950_o;
  wire n953_o;
  wire n956_o;
  wire n959_o;
  wire n962_o;
  wire n965_o;
  wire n968_o;
  wire n971_o;
  wire n974_o;
  wire n977_o;
  wire n980_o;
  wire n983_o;
  wire n986_o;
  wire n989_o;
  wire n992_o;
  wire n995_o;
  wire n998_o;
  wire n1001_o;
  wire n1004_o;
  wire n1007_o;
  wire n1010_o;
  wire n1013_o;
  wire n1016_o;
  wire n1019_o;
  wire n1022_o;
  wire n1025_o;
  wire n1028_o;
  wire n1031_o;
  wire n1034_o;
  wire n1037_o;
  wire n1040_o;
  wire n1043_o;
  wire n1046_o;
  wire n1049_o;
  wire n1052_o;
  wire n1055_o;
  wire n1058_o;
  wire n1061_o;
  wire n1064_o;
  wire n1067_o;
  wire n1070_o;
  wire n1073_o;
  wire n1076_o;
  wire n1079_o;
  wire n1082_o;
  wire n1085_o;
  wire n1088_o;
  wire n1091_o;
  wire n1094_o;
  wire n1097_o;
  wire n1100_o;
  wire n1103_o;
  wire n1106_o;
  wire n1109_o;
  wire n1112_o;
  wire n1115_o;
  wire n1118_o;
  wire n1121_o;
  wire n1124_o;
  wire n1127_o;
  wire n1130_o;
  wire n1133_o;
  wire n1136_o;
  wire n1139_o;
  wire n1142_o;
  wire n1145_o;
  wire n1148_o;
  wire n1151_o;
  wire n1154_o;
  wire n1157_o;
  wire n1160_o;
  wire n1163_o;
  wire n1166_o;
  wire n1169_o;
  wire n1172_o;
  wire n1175_o;
  wire n1178_o;
  wire n1181_o;
  wire n1184_o;
  wire n1187_o;
  wire n1190_o;
  wire n1193_o;
  wire n1196_o;
  wire n1199_o;
  wire n1202_o;
  wire n1205_o;
  wire n1208_o;
  wire n1211_o;
  wire n1214_o;
  wire n1217_o;
  wire n1220_o;
  wire n1223_o;
  wire n1226_o;
  wire n1229_o;
  wire n1232_o;
  wire n1235_o;
  wire n1238_o;
  wire n1241_o;
  wire n1244_o;
  wire n1247_o;
  wire n1250_o;
  wire n1253_o;
  wire n1256_o;
  wire n1259_o;
  wire n1262_o;
  wire n1265_o;
  wire n1268_o;
  wire n1271_o;
  wire n1274_o;
  wire n1277_o;
  wire n1280_o;
  wire n1283_o;
  wire n1286_o;
  wire n1289_o;
  wire n1292_o;
  wire n1295_o;
  wire n1298_o;
  wire n1301_o;
  wire n1304_o;
  wire n1307_o;
  wire n1310_o;
  wire n1313_o;
  wire n1316_o;
  wire n1319_o;
  wire n1322_o;
  wire n1325_o;
  wire n1328_o;
  wire n1331_o;
  wire n1334_o;
  wire n1337_o;
  wire n1340_o;
  wire n1343_o;
  wire n1346_o;
  wire n1349_o;
  wire n1352_o;
  wire n1355_o;
  wire n1358_o;
  wire n1361_o;
  wire n1364_o;
  wire n1367_o;
  wire n1370_o;
  wire n1373_o;
  wire n1376_o;
  wire n1379_o;
  wire n1382_o;
  wire n1385_o;
  wire n1388_o;
  wire n1391_o;
  wire n1394_o;
  wire n1397_o;
  wire n1400_o;
  wire n1403_o;
  wire n1406_o;
  wire n1409_o;
  wire n1412_o;
  wire n1415_o;
  wire n1418_o;
  wire n1421_o;
  wire n1424_o;
  wire n1427_o;
  wire n1430_o;
  wire n1433_o;
  wire n1436_o;
  wire n1439_o;
  wire n1442_o;
  wire n1445_o;
  wire n1448_o;
  wire n1451_o;
  wire n1454_o;
  wire n1457_o;
  wire n1460_o;
  wire n1463_o;
  wire n1466_o;
  wire n1469_o;
  wire n1472_o;
  wire n1475_o;
  wire n1478_o;
  wire n1481_o;
  wire n1484_o;
  wire n1487_o;
  wire n1490_o;
  wire n1493_o;
  wire n1496_o;
  wire n1499_o;
  wire n1502_o;
  wire n1505_o;
  wire n1508_o;
  wire n1511_o;
  wire n1514_o;
  wire n1517_o;
  wire n1520_o;
  wire n1523_o;
  wire n1526_o;
  wire n1529_o;
  wire n1532_o;
  wire n1535_o;
  wire n1538_o;
  wire n1541_o;
  wire n1544_o;
  wire n1547_o;
  wire n1550_o;
  wire n1553_o;
  wire n1556_o;
  wire n1559_o;
  wire n1562_o;
  wire n1565_o;
  wire n1568_o;
  wire n1571_o;
  wire n1574_o;
  wire n1577_o;
  wire n1580_o;
  wire n1583_o;
  wire n1586_o;
  wire n1589_o;
  wire n1592_o;
  wire n1595_o;
  wire n1598_o;
  wire n1601_o;
  wire n1604_o;
  wire n1607_o;
  wire n1610_o;
  wire n1613_o;
  wire n1616_o;
  wire n1619_o;
  wire n1622_o;
  wire n1625_o;
  wire n1628_o;
  wire n1631_o;
  wire n1634_o;
  wire n1637_o;
  wire n1640_o;
  wire n1643_o;
  wire n1646_o;
  wire n1649_o;
  wire n1652_o;
  wire n1655_o;
  wire n1658_o;
  wire n1661_o;
  wire n1664_o;
  wire n1667_o;
  wire n1670_o;
  wire n1673_o;
  wire n1676_o;
  wire n1679_o;
  wire n1682_o;
  wire n1685_o;
  wire n1688_o;
  wire n1691_o;
  wire n1694_o;
  wire n1697_o;
  wire n1700_o;
  wire n1703_o;
  wire n1706_o;
  wire n1709_o;
  wire n1712_o;
  wire n1715_o;
  wire n1718_o;
  wire n1721_o;
  wire n1724_o;
  wire n1727_o;
  wire n1730_o;
  wire n1733_o;
  wire n1736_o;
  wire n1739_o;
  wire n1742_o;
  wire n1745_o;
  wire n1748_o;
  wire n1751_o;
  wire n1754_o;
  wire n1757_o;
  wire n1760_o;
  wire n1763_o;
  wire n1766_o;
  wire n1769_o;
  wire n1772_o;
  wire n1775_o;
  wire n1778_o;
  wire n1781_o;
  wire n1784_o;
  wire n1787_o;
  wire n1790_o;
  wire n1793_o;
  wire n1796_o;
  wire n1799_o;
  wire n1802_o;
  wire n1805_o;
  wire n1808_o;
  wire n1811_o;
  wire n1814_o;
  wire n1817_o;
  wire n1820_o;
  wire n1823_o;
  wire n1826_o;
  wire n1829_o;
  wire n1832_o;
  wire n1835_o;
  wire n1838_o;
  wire n1841_o;
  wire n1844_o;
  wire n1847_o;
  wire n1850_o;
  wire n1853_o;
  wire n1856_o;
  wire n1859_o;
  wire n1862_o;
  wire n1865_o;
  wire n1868_o;
  wire n1871_o;
  wire n1874_o;
  wire n1877_o;
  wire n1880_o;
  wire n1883_o;
  wire n1886_o;
  wire n1889_o;
  wire n1892_o;
  wire n1895_o;
  wire n1898_o;
  wire n1901_o;
  wire n1904_o;
  wire n1907_o;
  wire n1910_o;
  wire n1913_o;
  wire n1916_o;
  wire n1919_o;
  wire n1922_o;
  wire n1925_o;
  wire n1928_o;
  wire n1931_o;
  wire n1934_o;
  wire n1937_o;
  wire n1940_o;
  wire n1943_o;
  wire n1946_o;
  wire n1949_o;
  wire n1952_o;
  wire n1955_o;
  wire n1958_o;
  wire n1961_o;
  wire n1964_o;
  wire n1967_o;
  wire n1970_o;
  wire n1973_o;
  wire n1976_o;
  wire n1979_o;
  wire n1982_o;
  wire n1985_o;
  wire n1988_o;
  wire n1991_o;
  wire n1994_o;
  wire n1997_o;
  wire n2000_o;
  wire n2003_o;
  wire n2006_o;
  wire n2009_o;
  wire n2012_o;
  wire n2015_o;
  wire n2018_o;
  wire n2021_o;
  wire n2024_o;
  wire n2027_o;
  wire n2030_o;
  wire n2033_o;
  wire n2036_o;
  wire n2039_o;
  wire n2042_o;
  wire [511:0] n2044_o;
  reg [2:0] n2045_o;
  assign y = y1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:28:8  */
  assign y0 = n2045_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:33:8  */
  assign y1 = y0; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:36:13  */
  assign n509_o = x == 9'b000000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:37:13  */
  assign n512_o = x == 9'b000000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:38:13  */
  assign n515_o = x == 9'b000000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:39:13  */
  assign n518_o = x == 9'b000000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:40:13  */
  assign n521_o = x == 9'b000000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:41:13  */
  assign n524_o = x == 9'b000000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:42:13  */
  assign n527_o = x == 9'b000000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:43:13  */
  assign n530_o = x == 9'b000000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:44:13  */
  assign n533_o = x == 9'b000001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:45:13  */
  assign n536_o = x == 9'b000001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:46:13  */
  assign n539_o = x == 9'b000001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:47:13  */
  assign n542_o = x == 9'b000001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:48:13  */
  assign n545_o = x == 9'b000001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:49:13  */
  assign n548_o = x == 9'b000001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:50:13  */
  assign n551_o = x == 9'b000001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:51:13  */
  assign n554_o = x == 9'b000001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:52:13  */
  assign n557_o = x == 9'b000010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:53:13  */
  assign n560_o = x == 9'b000010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:54:13  */
  assign n563_o = x == 9'b000010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:55:13  */
  assign n566_o = x == 9'b000010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:56:13  */
  assign n569_o = x == 9'b000010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:57:13  */
  assign n572_o = x == 9'b000010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:58:13  */
  assign n575_o = x == 9'b000010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:59:13  */
  assign n578_o = x == 9'b000010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:60:13  */
  assign n581_o = x == 9'b000011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:61:13  */
  assign n584_o = x == 9'b000011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:62:13  */
  assign n587_o = x == 9'b000011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:63:13  */
  assign n590_o = x == 9'b000011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:64:13  */
  assign n593_o = x == 9'b000011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:65:13  */
  assign n596_o = x == 9'b000011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:66:13  */
  assign n599_o = x == 9'b000011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:67:13  */
  assign n602_o = x == 9'b000011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:68:13  */
  assign n605_o = x == 9'b000100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:69:13  */
  assign n608_o = x == 9'b000100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:70:13  */
  assign n611_o = x == 9'b000100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:71:13  */
  assign n614_o = x == 9'b000100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:72:13  */
  assign n617_o = x == 9'b000100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:73:13  */
  assign n620_o = x == 9'b000100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:74:13  */
  assign n623_o = x == 9'b000100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:75:13  */
  assign n626_o = x == 9'b000100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:76:13  */
  assign n629_o = x == 9'b000101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:77:13  */
  assign n632_o = x == 9'b000101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:78:13  */
  assign n635_o = x == 9'b000101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:79:13  */
  assign n638_o = x == 9'b000101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:80:13  */
  assign n641_o = x == 9'b000101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:81:13  */
  assign n644_o = x == 9'b000101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:82:13  */
  assign n647_o = x == 9'b000101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:83:13  */
  assign n650_o = x == 9'b000101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:84:13  */
  assign n653_o = x == 9'b000110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:85:13  */
  assign n656_o = x == 9'b000110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:86:13  */
  assign n659_o = x == 9'b000110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:87:13  */
  assign n662_o = x == 9'b000110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:88:13  */
  assign n665_o = x == 9'b000110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:89:13  */
  assign n668_o = x == 9'b000110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:90:13  */
  assign n671_o = x == 9'b000110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:91:13  */
  assign n674_o = x == 9'b000110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:92:13  */
  assign n677_o = x == 9'b000111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:93:13  */
  assign n680_o = x == 9'b000111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:94:13  */
  assign n683_o = x == 9'b000111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:95:13  */
  assign n686_o = x == 9'b000111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:96:13  */
  assign n689_o = x == 9'b000111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:97:13  */
  assign n692_o = x == 9'b000111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:98:13  */
  assign n695_o = x == 9'b000111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:99:13  */
  assign n698_o = x == 9'b000111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:100:13  */
  assign n701_o = x == 9'b001000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:101:13  */
  assign n704_o = x == 9'b001000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:102:13  */
  assign n707_o = x == 9'b001000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:103:13  */
  assign n710_o = x == 9'b001000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:104:13  */
  assign n713_o = x == 9'b001000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:105:13  */
  assign n716_o = x == 9'b001000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:106:13  */
  assign n719_o = x == 9'b001000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:107:13  */
  assign n722_o = x == 9'b001000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:108:13  */
  assign n725_o = x == 9'b001001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:109:13  */
  assign n728_o = x == 9'b001001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:110:13  */
  assign n731_o = x == 9'b001001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:111:13  */
  assign n734_o = x == 9'b001001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:112:13  */
  assign n737_o = x == 9'b001001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:113:13  */
  assign n740_o = x == 9'b001001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:114:13  */
  assign n743_o = x == 9'b001001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:115:13  */
  assign n746_o = x == 9'b001001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:116:13  */
  assign n749_o = x == 9'b001010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:117:13  */
  assign n752_o = x == 9'b001010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:118:13  */
  assign n755_o = x == 9'b001010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:119:13  */
  assign n758_o = x == 9'b001010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:120:13  */
  assign n761_o = x == 9'b001010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:121:13  */
  assign n764_o = x == 9'b001010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:122:13  */
  assign n767_o = x == 9'b001010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:123:13  */
  assign n770_o = x == 9'b001010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:124:13  */
  assign n773_o = x == 9'b001011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:125:13  */
  assign n776_o = x == 9'b001011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:126:13  */
  assign n779_o = x == 9'b001011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:127:13  */
  assign n782_o = x == 9'b001011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:128:13  */
  assign n785_o = x == 9'b001011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:129:13  */
  assign n788_o = x == 9'b001011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:130:13  */
  assign n791_o = x == 9'b001011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:131:13  */
  assign n794_o = x == 9'b001011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:132:13  */
  assign n797_o = x == 9'b001100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:133:13  */
  assign n800_o = x == 9'b001100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:134:13  */
  assign n803_o = x == 9'b001100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:135:13  */
  assign n806_o = x == 9'b001100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:136:13  */
  assign n809_o = x == 9'b001100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:137:13  */
  assign n812_o = x == 9'b001100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:138:13  */
  assign n815_o = x == 9'b001100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:139:13  */
  assign n818_o = x == 9'b001100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:140:13  */
  assign n821_o = x == 9'b001101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:141:13  */
  assign n824_o = x == 9'b001101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:142:13  */
  assign n827_o = x == 9'b001101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:143:13  */
  assign n830_o = x == 9'b001101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:144:13  */
  assign n833_o = x == 9'b001101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:145:13  */
  assign n836_o = x == 9'b001101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:146:13  */
  assign n839_o = x == 9'b001101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:147:13  */
  assign n842_o = x == 9'b001101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:148:13  */
  assign n845_o = x == 9'b001110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:149:13  */
  assign n848_o = x == 9'b001110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:150:13  */
  assign n851_o = x == 9'b001110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:151:13  */
  assign n854_o = x == 9'b001110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:152:13  */
  assign n857_o = x == 9'b001110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:153:13  */
  assign n860_o = x == 9'b001110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:154:13  */
  assign n863_o = x == 9'b001110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:155:13  */
  assign n866_o = x == 9'b001110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:156:13  */
  assign n869_o = x == 9'b001111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:157:13  */
  assign n872_o = x == 9'b001111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:158:13  */
  assign n875_o = x == 9'b001111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:159:13  */
  assign n878_o = x == 9'b001111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:160:13  */
  assign n881_o = x == 9'b001111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:161:13  */
  assign n884_o = x == 9'b001111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:162:13  */
  assign n887_o = x == 9'b001111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:163:13  */
  assign n890_o = x == 9'b001111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:164:13  */
  assign n893_o = x == 9'b010000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:165:13  */
  assign n896_o = x == 9'b010000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:166:13  */
  assign n899_o = x == 9'b010000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:167:13  */
  assign n902_o = x == 9'b010000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:168:13  */
  assign n905_o = x == 9'b010000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:169:13  */
  assign n908_o = x == 9'b010000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:170:13  */
  assign n911_o = x == 9'b010000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:171:13  */
  assign n914_o = x == 9'b010000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:172:13  */
  assign n917_o = x == 9'b010001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:173:13  */
  assign n920_o = x == 9'b010001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:174:13  */
  assign n923_o = x == 9'b010001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:175:13  */
  assign n926_o = x == 9'b010001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:176:13  */
  assign n929_o = x == 9'b010001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:177:13  */
  assign n932_o = x == 9'b010001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:178:13  */
  assign n935_o = x == 9'b010001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:179:13  */
  assign n938_o = x == 9'b010001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:180:13  */
  assign n941_o = x == 9'b010010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:181:13  */
  assign n944_o = x == 9'b010010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:182:13  */
  assign n947_o = x == 9'b010010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:183:13  */
  assign n950_o = x == 9'b010010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:184:13  */
  assign n953_o = x == 9'b010010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:185:13  */
  assign n956_o = x == 9'b010010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:186:13  */
  assign n959_o = x == 9'b010010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:187:13  */
  assign n962_o = x == 9'b010010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:188:13  */
  assign n965_o = x == 9'b010011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:189:13  */
  assign n968_o = x == 9'b010011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:190:13  */
  assign n971_o = x == 9'b010011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:191:13  */
  assign n974_o = x == 9'b010011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:192:13  */
  assign n977_o = x == 9'b010011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:193:13  */
  assign n980_o = x == 9'b010011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:194:13  */
  assign n983_o = x == 9'b010011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:195:13  */
  assign n986_o = x == 9'b010011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:196:13  */
  assign n989_o = x == 9'b010100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:197:13  */
  assign n992_o = x == 9'b010100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:198:13  */
  assign n995_o = x == 9'b010100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:199:13  */
  assign n998_o = x == 9'b010100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:200:13  */
  assign n1001_o = x == 9'b010100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:201:13  */
  assign n1004_o = x == 9'b010100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:202:13  */
  assign n1007_o = x == 9'b010100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:203:13  */
  assign n1010_o = x == 9'b010100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:204:13  */
  assign n1013_o = x == 9'b010101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:205:13  */
  assign n1016_o = x == 9'b010101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:206:13  */
  assign n1019_o = x == 9'b010101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:207:13  */
  assign n1022_o = x == 9'b010101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:208:13  */
  assign n1025_o = x == 9'b010101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:209:13  */
  assign n1028_o = x == 9'b010101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:210:13  */
  assign n1031_o = x == 9'b010101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:211:13  */
  assign n1034_o = x == 9'b010101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:212:13  */
  assign n1037_o = x == 9'b010110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:213:13  */
  assign n1040_o = x == 9'b010110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:214:13  */
  assign n1043_o = x == 9'b010110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:215:13  */
  assign n1046_o = x == 9'b010110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:216:13  */
  assign n1049_o = x == 9'b010110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:217:13  */
  assign n1052_o = x == 9'b010110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:218:13  */
  assign n1055_o = x == 9'b010110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:219:13  */
  assign n1058_o = x == 9'b010110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:220:13  */
  assign n1061_o = x == 9'b010111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:221:13  */
  assign n1064_o = x == 9'b010111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:222:13  */
  assign n1067_o = x == 9'b010111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:223:13  */
  assign n1070_o = x == 9'b010111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:224:13  */
  assign n1073_o = x == 9'b010111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:225:13  */
  assign n1076_o = x == 9'b010111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:226:13  */
  assign n1079_o = x == 9'b010111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:227:13  */
  assign n1082_o = x == 9'b010111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:228:13  */
  assign n1085_o = x == 9'b011000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:229:13  */
  assign n1088_o = x == 9'b011000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:230:13  */
  assign n1091_o = x == 9'b011000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:231:13  */
  assign n1094_o = x == 9'b011000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:232:13  */
  assign n1097_o = x == 9'b011000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:233:13  */
  assign n1100_o = x == 9'b011000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:234:13  */
  assign n1103_o = x == 9'b011000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:235:13  */
  assign n1106_o = x == 9'b011000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:236:13  */
  assign n1109_o = x == 9'b011001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:237:13  */
  assign n1112_o = x == 9'b011001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:238:13  */
  assign n1115_o = x == 9'b011001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:239:13  */
  assign n1118_o = x == 9'b011001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:240:13  */
  assign n1121_o = x == 9'b011001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:241:13  */
  assign n1124_o = x == 9'b011001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:242:13  */
  assign n1127_o = x == 9'b011001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:243:13  */
  assign n1130_o = x == 9'b011001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:244:13  */
  assign n1133_o = x == 9'b011010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:245:13  */
  assign n1136_o = x == 9'b011010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:246:13  */
  assign n1139_o = x == 9'b011010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:247:13  */
  assign n1142_o = x == 9'b011010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:248:13  */
  assign n1145_o = x == 9'b011010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:249:13  */
  assign n1148_o = x == 9'b011010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:250:13  */
  assign n1151_o = x == 9'b011010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:251:13  */
  assign n1154_o = x == 9'b011010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:252:13  */
  assign n1157_o = x == 9'b011011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:253:13  */
  assign n1160_o = x == 9'b011011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:254:13  */
  assign n1163_o = x == 9'b011011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:255:13  */
  assign n1166_o = x == 9'b011011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:256:13  */
  assign n1169_o = x == 9'b011011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:257:13  */
  assign n1172_o = x == 9'b011011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:258:13  */
  assign n1175_o = x == 9'b011011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:259:13  */
  assign n1178_o = x == 9'b011011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:260:13  */
  assign n1181_o = x == 9'b011100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:261:13  */
  assign n1184_o = x == 9'b011100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:262:13  */
  assign n1187_o = x == 9'b011100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:263:13  */
  assign n1190_o = x == 9'b011100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:264:13  */
  assign n1193_o = x == 9'b011100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:265:13  */
  assign n1196_o = x == 9'b011100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:266:13  */
  assign n1199_o = x == 9'b011100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:267:13  */
  assign n1202_o = x == 9'b011100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:268:13  */
  assign n1205_o = x == 9'b011101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:269:13  */
  assign n1208_o = x == 9'b011101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:270:13  */
  assign n1211_o = x == 9'b011101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:271:13  */
  assign n1214_o = x == 9'b011101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:272:13  */
  assign n1217_o = x == 9'b011101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:273:13  */
  assign n1220_o = x == 9'b011101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:274:13  */
  assign n1223_o = x == 9'b011101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:275:13  */
  assign n1226_o = x == 9'b011101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:276:13  */
  assign n1229_o = x == 9'b011110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:277:13  */
  assign n1232_o = x == 9'b011110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:278:13  */
  assign n1235_o = x == 9'b011110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:279:13  */
  assign n1238_o = x == 9'b011110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:280:13  */
  assign n1241_o = x == 9'b011110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:281:13  */
  assign n1244_o = x == 9'b011110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:282:13  */
  assign n1247_o = x == 9'b011110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:283:13  */
  assign n1250_o = x == 9'b011110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:284:13  */
  assign n1253_o = x == 9'b011111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:285:13  */
  assign n1256_o = x == 9'b011111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:286:13  */
  assign n1259_o = x == 9'b011111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:287:13  */
  assign n1262_o = x == 9'b011111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:288:13  */
  assign n1265_o = x == 9'b011111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:289:13  */
  assign n1268_o = x == 9'b011111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:290:13  */
  assign n1271_o = x == 9'b011111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:291:13  */
  assign n1274_o = x == 9'b011111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:292:13  */
  assign n1277_o = x == 9'b100000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:293:13  */
  assign n1280_o = x == 9'b100000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:294:13  */
  assign n1283_o = x == 9'b100000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:295:13  */
  assign n1286_o = x == 9'b100000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:296:13  */
  assign n1289_o = x == 9'b100000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:297:13  */
  assign n1292_o = x == 9'b100000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:298:13  */
  assign n1295_o = x == 9'b100000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:299:13  */
  assign n1298_o = x == 9'b100000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:300:13  */
  assign n1301_o = x == 9'b100001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:301:13  */
  assign n1304_o = x == 9'b100001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:302:13  */
  assign n1307_o = x == 9'b100001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:303:13  */
  assign n1310_o = x == 9'b100001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:304:13  */
  assign n1313_o = x == 9'b100001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:305:13  */
  assign n1316_o = x == 9'b100001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:306:13  */
  assign n1319_o = x == 9'b100001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:307:13  */
  assign n1322_o = x == 9'b100001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:308:13  */
  assign n1325_o = x == 9'b100010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:309:13  */
  assign n1328_o = x == 9'b100010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:310:13  */
  assign n1331_o = x == 9'b100010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:311:13  */
  assign n1334_o = x == 9'b100010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:312:13  */
  assign n1337_o = x == 9'b100010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:313:13  */
  assign n1340_o = x == 9'b100010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:314:13  */
  assign n1343_o = x == 9'b100010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:315:13  */
  assign n1346_o = x == 9'b100010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:316:13  */
  assign n1349_o = x == 9'b100011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:317:13  */
  assign n1352_o = x == 9'b100011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:318:13  */
  assign n1355_o = x == 9'b100011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:319:13  */
  assign n1358_o = x == 9'b100011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:320:13  */
  assign n1361_o = x == 9'b100011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:321:13  */
  assign n1364_o = x == 9'b100011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:322:13  */
  assign n1367_o = x == 9'b100011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:323:13  */
  assign n1370_o = x == 9'b100011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:324:13  */
  assign n1373_o = x == 9'b100100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:325:13  */
  assign n1376_o = x == 9'b100100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:326:13  */
  assign n1379_o = x == 9'b100100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:327:13  */
  assign n1382_o = x == 9'b100100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:328:13  */
  assign n1385_o = x == 9'b100100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:329:13  */
  assign n1388_o = x == 9'b100100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:330:13  */
  assign n1391_o = x == 9'b100100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:331:13  */
  assign n1394_o = x == 9'b100100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:332:13  */
  assign n1397_o = x == 9'b100101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:333:13  */
  assign n1400_o = x == 9'b100101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:334:13  */
  assign n1403_o = x == 9'b100101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:335:13  */
  assign n1406_o = x == 9'b100101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:336:13  */
  assign n1409_o = x == 9'b100101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:337:13  */
  assign n1412_o = x == 9'b100101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:338:13  */
  assign n1415_o = x == 9'b100101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:339:13  */
  assign n1418_o = x == 9'b100101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:340:13  */
  assign n1421_o = x == 9'b100110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:341:13  */
  assign n1424_o = x == 9'b100110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:342:13  */
  assign n1427_o = x == 9'b100110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:343:13  */
  assign n1430_o = x == 9'b100110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:344:13  */
  assign n1433_o = x == 9'b100110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:345:13  */
  assign n1436_o = x == 9'b100110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:346:13  */
  assign n1439_o = x == 9'b100110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:347:13  */
  assign n1442_o = x == 9'b100110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:348:13  */
  assign n1445_o = x == 9'b100111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:349:13  */
  assign n1448_o = x == 9'b100111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:350:13  */
  assign n1451_o = x == 9'b100111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:351:13  */
  assign n1454_o = x == 9'b100111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:352:13  */
  assign n1457_o = x == 9'b100111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:353:13  */
  assign n1460_o = x == 9'b100111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:354:13  */
  assign n1463_o = x == 9'b100111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:355:13  */
  assign n1466_o = x == 9'b100111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:356:13  */
  assign n1469_o = x == 9'b101000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:357:13  */
  assign n1472_o = x == 9'b101000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:358:13  */
  assign n1475_o = x == 9'b101000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:359:13  */
  assign n1478_o = x == 9'b101000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:360:13  */
  assign n1481_o = x == 9'b101000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:361:13  */
  assign n1484_o = x == 9'b101000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:362:13  */
  assign n1487_o = x == 9'b101000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:363:13  */
  assign n1490_o = x == 9'b101000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:364:13  */
  assign n1493_o = x == 9'b101001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:365:13  */
  assign n1496_o = x == 9'b101001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:366:13  */
  assign n1499_o = x == 9'b101001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:367:13  */
  assign n1502_o = x == 9'b101001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:368:13  */
  assign n1505_o = x == 9'b101001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:369:13  */
  assign n1508_o = x == 9'b101001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:370:13  */
  assign n1511_o = x == 9'b101001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:371:13  */
  assign n1514_o = x == 9'b101001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:372:13  */
  assign n1517_o = x == 9'b101010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:373:13  */
  assign n1520_o = x == 9'b101010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:374:13  */
  assign n1523_o = x == 9'b101010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:375:13  */
  assign n1526_o = x == 9'b101010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:376:13  */
  assign n1529_o = x == 9'b101010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:377:13  */
  assign n1532_o = x == 9'b101010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:378:13  */
  assign n1535_o = x == 9'b101010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:379:13  */
  assign n1538_o = x == 9'b101010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:380:13  */
  assign n1541_o = x == 9'b101011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:381:13  */
  assign n1544_o = x == 9'b101011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:382:13  */
  assign n1547_o = x == 9'b101011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:383:13  */
  assign n1550_o = x == 9'b101011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:384:13  */
  assign n1553_o = x == 9'b101011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:385:13  */
  assign n1556_o = x == 9'b101011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:386:13  */
  assign n1559_o = x == 9'b101011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:387:13  */
  assign n1562_o = x == 9'b101011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:388:13  */
  assign n1565_o = x == 9'b101100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:389:13  */
  assign n1568_o = x == 9'b101100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:390:13  */
  assign n1571_o = x == 9'b101100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:391:13  */
  assign n1574_o = x == 9'b101100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:392:13  */
  assign n1577_o = x == 9'b101100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:393:13  */
  assign n1580_o = x == 9'b101100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:394:13  */
  assign n1583_o = x == 9'b101100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:395:13  */
  assign n1586_o = x == 9'b101100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:396:13  */
  assign n1589_o = x == 9'b101101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:397:13  */
  assign n1592_o = x == 9'b101101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:398:13  */
  assign n1595_o = x == 9'b101101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:399:13  */
  assign n1598_o = x == 9'b101101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:400:13  */
  assign n1601_o = x == 9'b101101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:401:13  */
  assign n1604_o = x == 9'b101101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:402:13  */
  assign n1607_o = x == 9'b101101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:403:13  */
  assign n1610_o = x == 9'b101101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:404:13  */
  assign n1613_o = x == 9'b101110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:405:13  */
  assign n1616_o = x == 9'b101110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:406:13  */
  assign n1619_o = x == 9'b101110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:407:13  */
  assign n1622_o = x == 9'b101110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:408:13  */
  assign n1625_o = x == 9'b101110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:409:13  */
  assign n1628_o = x == 9'b101110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:410:13  */
  assign n1631_o = x == 9'b101110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:411:13  */
  assign n1634_o = x == 9'b101110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:412:13  */
  assign n1637_o = x == 9'b101111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:413:13  */
  assign n1640_o = x == 9'b101111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:414:13  */
  assign n1643_o = x == 9'b101111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:415:13  */
  assign n1646_o = x == 9'b101111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:416:13  */
  assign n1649_o = x == 9'b101111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:417:13  */
  assign n1652_o = x == 9'b101111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:418:13  */
  assign n1655_o = x == 9'b101111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:419:13  */
  assign n1658_o = x == 9'b101111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:420:13  */
  assign n1661_o = x == 9'b110000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:421:13  */
  assign n1664_o = x == 9'b110000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:422:13  */
  assign n1667_o = x == 9'b110000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:423:13  */
  assign n1670_o = x == 9'b110000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:424:13  */
  assign n1673_o = x == 9'b110000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:425:13  */
  assign n1676_o = x == 9'b110000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:426:13  */
  assign n1679_o = x == 9'b110000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:427:13  */
  assign n1682_o = x == 9'b110000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:428:13  */
  assign n1685_o = x == 9'b110001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:429:13  */
  assign n1688_o = x == 9'b110001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:430:13  */
  assign n1691_o = x == 9'b110001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:431:13  */
  assign n1694_o = x == 9'b110001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:432:13  */
  assign n1697_o = x == 9'b110001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:433:13  */
  assign n1700_o = x == 9'b110001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:434:13  */
  assign n1703_o = x == 9'b110001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:435:13  */
  assign n1706_o = x == 9'b110001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:436:13  */
  assign n1709_o = x == 9'b110010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:437:13  */
  assign n1712_o = x == 9'b110010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:438:13  */
  assign n1715_o = x == 9'b110010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:439:13  */
  assign n1718_o = x == 9'b110010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:440:13  */
  assign n1721_o = x == 9'b110010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:441:13  */
  assign n1724_o = x == 9'b110010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:442:13  */
  assign n1727_o = x == 9'b110010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:443:13  */
  assign n1730_o = x == 9'b110010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:444:13  */
  assign n1733_o = x == 9'b110011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:445:13  */
  assign n1736_o = x == 9'b110011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:446:13  */
  assign n1739_o = x == 9'b110011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:447:13  */
  assign n1742_o = x == 9'b110011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:448:13  */
  assign n1745_o = x == 9'b110011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:449:13  */
  assign n1748_o = x == 9'b110011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:450:13  */
  assign n1751_o = x == 9'b110011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:451:13  */
  assign n1754_o = x == 9'b110011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:452:13  */
  assign n1757_o = x == 9'b110100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:453:13  */
  assign n1760_o = x == 9'b110100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:454:13  */
  assign n1763_o = x == 9'b110100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:455:13  */
  assign n1766_o = x == 9'b110100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:456:13  */
  assign n1769_o = x == 9'b110100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:457:13  */
  assign n1772_o = x == 9'b110100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:458:13  */
  assign n1775_o = x == 9'b110100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:459:13  */
  assign n1778_o = x == 9'b110100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:460:13  */
  assign n1781_o = x == 9'b110101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:461:13  */
  assign n1784_o = x == 9'b110101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:462:13  */
  assign n1787_o = x == 9'b110101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:463:13  */
  assign n1790_o = x == 9'b110101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:464:13  */
  assign n1793_o = x == 9'b110101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:465:13  */
  assign n1796_o = x == 9'b110101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:466:13  */
  assign n1799_o = x == 9'b110101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:467:13  */
  assign n1802_o = x == 9'b110101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:468:13  */
  assign n1805_o = x == 9'b110110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:469:13  */
  assign n1808_o = x == 9'b110110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:470:13  */
  assign n1811_o = x == 9'b110110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:471:13  */
  assign n1814_o = x == 9'b110110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:472:13  */
  assign n1817_o = x == 9'b110110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:473:13  */
  assign n1820_o = x == 9'b110110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:474:13  */
  assign n1823_o = x == 9'b110110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:475:13  */
  assign n1826_o = x == 9'b110110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:476:13  */
  assign n1829_o = x == 9'b110111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:477:13  */
  assign n1832_o = x == 9'b110111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:478:13  */
  assign n1835_o = x == 9'b110111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:479:13  */
  assign n1838_o = x == 9'b110111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:480:13  */
  assign n1841_o = x == 9'b110111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:481:13  */
  assign n1844_o = x == 9'b110111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:482:13  */
  assign n1847_o = x == 9'b110111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:483:13  */
  assign n1850_o = x == 9'b110111111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:484:13  */
  assign n1853_o = x == 9'b111000000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:485:13  */
  assign n1856_o = x == 9'b111000001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:486:13  */
  assign n1859_o = x == 9'b111000010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:487:13  */
  assign n1862_o = x == 9'b111000011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:488:13  */
  assign n1865_o = x == 9'b111000100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:489:13  */
  assign n1868_o = x == 9'b111000101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:490:13  */
  assign n1871_o = x == 9'b111000110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:491:13  */
  assign n1874_o = x == 9'b111000111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:492:13  */
  assign n1877_o = x == 9'b111001000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:493:13  */
  assign n1880_o = x == 9'b111001001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:494:13  */
  assign n1883_o = x == 9'b111001010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:495:13  */
  assign n1886_o = x == 9'b111001011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:496:13  */
  assign n1889_o = x == 9'b111001100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:497:13  */
  assign n1892_o = x == 9'b111001101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:498:13  */
  assign n1895_o = x == 9'b111001110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:499:13  */
  assign n1898_o = x == 9'b111001111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:500:13  */
  assign n1901_o = x == 9'b111010000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:501:13  */
  assign n1904_o = x == 9'b111010001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:502:13  */
  assign n1907_o = x == 9'b111010010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:503:13  */
  assign n1910_o = x == 9'b111010011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:504:13  */
  assign n1913_o = x == 9'b111010100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:505:13  */
  assign n1916_o = x == 9'b111010101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:506:13  */
  assign n1919_o = x == 9'b111010110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:507:13  */
  assign n1922_o = x == 9'b111010111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:508:13  */
  assign n1925_o = x == 9'b111011000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:509:13  */
  assign n1928_o = x == 9'b111011001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:510:13  */
  assign n1931_o = x == 9'b111011010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:511:13  */
  assign n1934_o = x == 9'b111011011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:512:13  */
  assign n1937_o = x == 9'b111011100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:513:13  */
  assign n1940_o = x == 9'b111011101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:514:13  */
  assign n1943_o = x == 9'b111011110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:515:13  */
  assign n1946_o = x == 9'b111011111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:516:13  */
  assign n1949_o = x == 9'b111100000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:517:13  */
  assign n1952_o = x == 9'b111100001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:518:13  */
  assign n1955_o = x == 9'b111100010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:519:13  */
  assign n1958_o = x == 9'b111100011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:520:13  */
  assign n1961_o = x == 9'b111100100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:521:13  */
  assign n1964_o = x == 9'b111100101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:522:13  */
  assign n1967_o = x == 9'b111100110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:523:13  */
  assign n1970_o = x == 9'b111100111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:524:13  */
  assign n1973_o = x == 9'b111101000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:525:13  */
  assign n1976_o = x == 9'b111101001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:526:13  */
  assign n1979_o = x == 9'b111101010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:527:13  */
  assign n1982_o = x == 9'b111101011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:528:13  */
  assign n1985_o = x == 9'b111101100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:529:13  */
  assign n1988_o = x == 9'b111101101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:530:13  */
  assign n1991_o = x == 9'b111101110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:531:13  */
  assign n1994_o = x == 9'b111101111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:532:13  */
  assign n1997_o = x == 9'b111110000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:533:13  */
  assign n2000_o = x == 9'b111110001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:534:13  */
  assign n2003_o = x == 9'b111110010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:535:13  */
  assign n2006_o = x == 9'b111110011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:536:13  */
  assign n2009_o = x == 9'b111110100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:537:13  */
  assign n2012_o = x == 9'b111110101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:538:13  */
  assign n2015_o = x == 9'b111110110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:539:13  */
  assign n2018_o = x == 9'b111110111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:540:13  */
  assign n2021_o = x == 9'b111111000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:541:13  */
  assign n2024_o = x == 9'b111111001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:542:13  */
  assign n2027_o = x == 9'b111111010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:543:13  */
  assign n2030_o = x == 9'b111111011;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:544:13  */
  assign n2033_o = x == 9'b111111100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:545:13  */
  assign n2036_o = x == 9'b111111101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:546:13  */
  assign n2039_o = x == 9'b111111110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:547:13  */
  assign n2042_o = x == 9'b111111111;
  assign n2044_o = {n2042_o, n2039_o, n2036_o, n2033_o, n2030_o, n2027_o, n2024_o, n2021_o, n2018_o, n2015_o, n2012_o, n2009_o, n2006_o, n2003_o, n2000_o, n1997_o, n1994_o, n1991_o, n1988_o, n1985_o, n1982_o, n1979_o, n1976_o, n1973_o, n1970_o, n1967_o, n1964_o, n1961_o, n1958_o, n1955_o, n1952_o, n1949_o, n1946_o, n1943_o, n1940_o, n1937_o, n1934_o, n1931_o, n1928_o, n1925_o, n1922_o, n1919_o, n1916_o, n1913_o, n1910_o, n1907_o, n1904_o, n1901_o, n1898_o, n1895_o, n1892_o, n1889_o, n1886_o, n1883_o, n1880_o, n1877_o, n1874_o, n1871_o, n1868_o, n1865_o, n1862_o, n1859_o, n1856_o, n1853_o, n1850_o, n1847_o, n1844_o, n1841_o, n1838_o, n1835_o, n1832_o, n1829_o, n1826_o, n1823_o, n1820_o, n1817_o, n1814_o, n1811_o, n1808_o, n1805_o, n1802_o, n1799_o, n1796_o, n1793_o, n1790_o, n1787_o, n1784_o, n1781_o, n1778_o, n1775_o, n1772_o, n1769_o, n1766_o, n1763_o, n1760_o, n1757_o, n1754_o, n1751_o, n1748_o, n1745_o, n1742_o, n1739_o, n1736_o, n1733_o, n1730_o, n1727_o, n1724_o, n1721_o, n1718_o, n1715_o, n1712_o, n1709_o, n1706_o, n1703_o, n1700_o, n1697_o, n1694_o, n1691_o, n1688_o, n1685_o, n1682_o, n1679_o, n1676_o, n1673_o, n1670_o, n1667_o, n1664_o, n1661_o, n1658_o, n1655_o, n1652_o, n1649_o, n1646_o, n1643_o, n1640_o, n1637_o, n1634_o, n1631_o, n1628_o, n1625_o, n1622_o, n1619_o, n1616_o, n1613_o, n1610_o, n1607_o, n1604_o, n1601_o, n1598_o, n1595_o, n1592_o, n1589_o, n1586_o, n1583_o, n1580_o, n1577_o, n1574_o, n1571_o, n1568_o, n1565_o, n1562_o, n1559_o, n1556_o, n1553_o, n1550_o, n1547_o, n1544_o, n1541_o, n1538_o, n1535_o, n1532_o, n1529_o, n1526_o, n1523_o, n1520_o, n1517_o, n1514_o, n1511_o, n1508_o, n1505_o, n1502_o, n1499_o, n1496_o, n1493_o, n1490_o, n1487_o, n1484_o, n1481_o, n1478_o, n1475_o, n1472_o, n1469_o, n1466_o, n1463_o, n1460_o, n1457_o, n1454_o, n1451_o, n1448_o, n1445_o, n1442_o, n1439_o, n1436_o, n1433_o, n1430_o, n1427_o, n1424_o, n1421_o, n1418_o, n1415_o, n1412_o, n1409_o, n1406_o, n1403_o, n1400_o, n1397_o, n1394_o, n1391_o, n1388_o, n1385_o, n1382_o, n1379_o, n1376_o, n1373_o, n1370_o, n1367_o, n1364_o, n1361_o, n1358_o, n1355_o, n1352_o, n1349_o, n1346_o, n1343_o, n1340_o, n1337_o, n1334_o, n1331_o, n1328_o, n1325_o, n1322_o, n1319_o, n1316_o, n1313_o, n1310_o, n1307_o, n1304_o, n1301_o, n1298_o, n1295_o, n1292_o, n1289_o, n1286_o, n1283_o, n1280_o, n1277_o, n1274_o, n1271_o, n1268_o, n1265_o, n1262_o, n1259_o, n1256_o, n1253_o, n1250_o, n1247_o, n1244_o, n1241_o, n1238_o, n1235_o, n1232_o, n1229_o, n1226_o, n1223_o, n1220_o, n1217_o, n1214_o, n1211_o, n1208_o, n1205_o, n1202_o, n1199_o, n1196_o, n1193_o, n1190_o, n1187_o, n1184_o, n1181_o, n1178_o, n1175_o, n1172_o, n1169_o, n1166_o, n1163_o, n1160_o, n1157_o, n1154_o, n1151_o, n1148_o, n1145_o, n1142_o, n1139_o, n1136_o, n1133_o, n1130_o, n1127_o, n1124_o, n1121_o, n1118_o, n1115_o, n1112_o, n1109_o, n1106_o, n1103_o, n1100_o, n1097_o, n1094_o, n1091_o, n1088_o, n1085_o, n1082_o, n1079_o, n1076_o, n1073_o, n1070_o, n1067_o, n1064_o, n1061_o, n1058_o, n1055_o, n1052_o, n1049_o, n1046_o, n1043_o, n1040_o, n1037_o, n1034_o, n1031_o, n1028_o, n1025_o, n1022_o, n1019_o, n1016_o, n1013_o, n1010_o, n1007_o, n1004_o, n1001_o, n998_o, n995_o, n992_o, n989_o, n986_o, n983_o, n980_o, n977_o, n974_o, n971_o, n968_o, n965_o, n962_o, n959_o, n956_o, n953_o, n950_o, n947_o, n944_o, n941_o, n938_o, n935_o, n932_o, n929_o, n926_o, n923_o, n920_o, n917_o, n914_o, n911_o, n908_o, n905_o, n902_o, n899_o, n896_o, n893_o, n890_o, n887_o, n884_o, n881_o, n878_o, n875_o, n872_o, n869_o, n866_o, n863_o, n860_o, n857_o, n854_o, n851_o, n848_o, n845_o, n842_o, n839_o, n836_o, n833_o, n830_o, n827_o, n824_o, n821_o, n818_o, n815_o, n812_o, n809_o, n806_o, n803_o, n800_o, n797_o, n794_o, n791_o, n788_o, n785_o, n782_o, n779_o, n776_o, n773_o, n770_o, n767_o, n764_o, n761_o, n758_o, n755_o, n752_o, n749_o, n746_o, n743_o, n740_o, n737_o, n734_o, n731_o, n728_o, n725_o, n722_o, n719_o, n716_o, n713_o, n710_o, n707_o, n704_o, n701_o, n698_o, n695_o, n692_o, n689_o, n686_o, n683_o, n680_o, n677_o, n674_o, n671_o, n668_o, n665_o, n662_o, n659_o, n656_o, n653_o, n650_o, n647_o, n644_o, n641_o, n638_o, n635_o, n632_o, n629_o, n626_o, n623_o, n620_o, n617_o, n614_o, n611_o, n608_o, n605_o, n602_o, n599_o, n596_o, n593_o, n590_o, n587_o, n584_o, n581_o, n578_o, n575_o, n572_o, n569_o, n566_o, n563_o, n560_o, n557_o, n554_o, n551_o, n548_o, n545_o, n542_o, n539_o, n536_o, n533_o, n530_o, n527_o, n524_o, n521_o, n518_o, n515_o, n512_o, n509_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:35:4  */
  always @*
    case (n2044_o)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2045_o = 3'b010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2045_o = 3'b001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2045_o = 3'b000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2045_o = 3'b000;
      default: n2045_o = 3'bXXX;
    endcase
endmodule

module fdiv #(parameter ID = 1)
  (input wire clk,
   input wire [16:0] X,
   input wire [16:0] Y,
   output wire [16:0] R);
  wire [10:0] fx;
  wire [10:0] fy;
  wire [5:0] expr0;
  wire [5:0] expr0_d1;
  wire [5:0] expr0_d2;
  wire [5:0] expr0_d3;
  wire [5:0] expr0_d4;
  wire [5:0] expr0_d5;
  wire [5:0] expr0_d6;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire [3:0] exnxy;
  wire [1:0] exnr0;
  wire [1:0] exnr0_d1;
  wire [1:0] exnr0_d2;
  wire [1:0] exnr0_d3;
  wire [1:0] exnr0_d4;
  wire [1:0] exnr0_d5;
  wire [1:0] exnr0_d6;
  wire [10:0] d;
  wire [10:0] d_d1;
  wire [10:0] d_d2;
  wire [10:0] d_d3;
  wire [10:0] d_d4;
  wire [10:0] d_d5;
  wire [11:0] psx;
  wire [13:0] betaw7;
  wire [8:0] sel7;
  wire [2:0] q7;
  wire [2:0] q7_copy5;
  wire [13:0] absq7d;
  wire [13:0] w6;
  wire [13:0] betaw6;
  wire [13:0] betaw6_d1;
  wire [8:0] sel6;
  wire [2:0] q6;
  wire [2:0] q6_copy6;
  wire [2:0] q6_copy6_d1;
  wire [13:0] absq6d;
  wire [13:0] w5;
  wire [13:0] betaw5;
  wire [13:0] betaw5_d1;
  wire [8:0] sel5;
  wire [2:0] q5;
  wire [2:0] q5_copy7;
  wire [2:0] q5_copy7_d1;
  wire [13:0] absq5d;
  wire [13:0] w4;
  wire [13:0] betaw4;
  wire [13:0] betaw4_d1;
  wire [8:0] sel4;
  wire [2:0] q4;
  wire [2:0] q4_d1;
  wire [2:0] q4_copy8;
  wire [13:0] absq4d;
  wire [13:0] absq4d_d1;
  wire [13:0] w3;
  wire [13:0] betaw3;
  wire [13:0] betaw3_d1;
  wire [8:0] sel3;
  wire [2:0] q3;
  wire [2:0] q3_d1;
  wire [2:0] q3_copy9;
  wire [13:0] absq3d;
  wire [13:0] absq3d_d1;
  wire [13:0] w2;
  wire [13:0] betaw2;
  wire [8:0] sel2;
  wire [2:0] q2;
  wire [2:0] q2_copy10;
  wire [13:0] absq2d;
  wire [13:0] w1;
  wire [13:0] betaw1;
  wire [13:0] betaw1_d1;
  wire [8:0] sel1;
  wire [2:0] q1;
  wire [2:0] q1_copy11;
  wire [2:0] q1_copy11_d1;
  wire [13:0] absq1d;
  wire [13:0] w0;
  wire [11:0] wfinal;
  wire qm0;
  wire [1:0] qp7;
  wire [1:0] qp7_d1;
  wire [1:0] qp7_d2;
  wire [1:0] qp7_d3;
  wire [1:0] qp7_d4;
  wire [1:0] qp7_d5;
  wire [1:0] qm7;
  wire [1:0] qm7_d1;
  wire [1:0] qm7_d2;
  wire [1:0] qm7_d3;
  wire [1:0] qm7_d4;
  wire [1:0] qm7_d5;
  wire [1:0] qp6;
  wire [1:0] qp6_d1;
  wire [1:0] qp6_d2;
  wire [1:0] qp6_d3;
  wire [1:0] qp6_d4;
  wire [1:0] qm6;
  wire [1:0] qm6_d1;
  wire [1:0] qm6_d2;
  wire [1:0] qm6_d3;
  wire [1:0] qm6_d4;
  wire [1:0] qp5;
  wire [1:0] qp5_d1;
  wire [1:0] qp5_d2;
  wire [1:0] qp5_d3;
  wire [1:0] qm5;
  wire [1:0] qm5_d1;
  wire [1:0] qm5_d2;
  wire [1:0] qm5_d3;
  wire [1:0] qp4;
  wire [1:0] qp4_d1;
  wire [1:0] qp4_d2;
  wire [1:0] qp4_d3;
  wire [1:0] qm4;
  wire [1:0] qm4_d1;
  wire [1:0] qm4_d2;
  wire [1:0] qm4_d3;
  wire [1:0] qp3;
  wire [1:0] qp3_d1;
  wire [1:0] qp3_d2;
  wire [1:0] qm3;
  wire [1:0] qm3_d1;
  wire [1:0] qm3_d2;
  wire [1:0] qp2;
  wire [1:0] qp2_d1;
  wire [1:0] qm2;
  wire [1:0] qm2_d1;
  wire [1:0] qp1;
  wire [1:0] qm1;
  wire [13:0] qp;
  wire [13:0] qm;
  wire [13:0] quotient;
  wire [13:0] quotient_d1;
  wire [12:0] mr;
  wire [10:0] frnorm;
  wire round;
  wire [5:0] expr1;
  wire [15:0] expfrac;
  wire [15:0] expfracr;
  wire [1:0] exnr;
  wire [1:0] exnrfinal;
  wire [9:0] n77_o;
  wire [10:0] n79_o;
  wire [9:0] n80_o;
  wire [10:0] n82_o;
  wire [3:0] n83_o;
  wire [5:0] n85_o;
  wire [3:0] n86_o;
  wire [5:0] n88_o;
  wire [5:0] n89_o;
  wire n90_o;
  wire n91_o;
  wire n92_o;
  wire [1:0] n93_o;
  wire [1:0] n94_o;
  wire [3:0] n95_o;
  wire n98_o;
  wire n101_o;
  wire n103_o;
  wire n104_o;
  wire n106_o;
  wire n107_o;
  wire n110_o;
  wire n112_o;
  wire n113_o;
  wire n115_o;
  wire n116_o;
  wire [2:0] n118_o;
  reg [1:0] n119_o;
  wire [11:0] n121_o;
  wire [13:0] n123_o;
  wire [5:0] n124_o;
  wire [2:0] n125_o;
  wire [8:0] n126_o;
  wire [2:0] selfunctiontable7_n127;
  wire [2:0] selfunctiontable7_y;
  wire [13:0] n131_o;
  wire n133_o;
  wire n135_o;
  wire n136_o;
  wire [12:0] n138_o;
  wire [13:0] n140_o;
  wire n142_o;
  wire n144_o;
  wire n145_o;
  wire [1:0] n147_o;
  reg [13:0] n148_o;
  wire n149_o;
  wire [13:0] n150_o;
  wire n152_o;
  wire [13:0] n153_o;
  reg [13:0] n154_o;
  wire [11:0] n155_o;
  wire [13:0] n157_o;
  wire [5:0] n158_o;
  wire [2:0] n159_o;
  wire [8:0] n160_o;
  wire [2:0] selfunctiontable6_n161;
  wire [2:0] selfunctiontable6_y;
  wire [13:0] n165_o;
  wire n167_o;
  wire n169_o;
  wire n170_o;
  wire [12:0] n172_o;
  wire [13:0] n174_o;
  wire n176_o;
  wire n178_o;
  wire n179_o;
  wire [1:0] n181_o;
  reg [13:0] n182_o;
  wire n183_o;
  wire [13:0] n184_o;
  wire n186_o;
  wire [13:0] n187_o;
  reg [13:0] n188_o;
  wire [11:0] n189_o;
  wire [13:0] n191_o;
  wire [5:0] n192_o;
  wire [2:0] n193_o;
  wire [8:0] n194_o;
  wire [2:0] selfunctiontable5_n195;
  wire [2:0] selfunctiontable5_y;
  wire [13:0] n199_o;
  wire n201_o;
  wire n203_o;
  wire n204_o;
  wire [12:0] n206_o;
  wire [13:0] n208_o;
  wire n210_o;
  wire n212_o;
  wire n213_o;
  wire [1:0] n215_o;
  reg [13:0] n216_o;
  wire n217_o;
  wire [13:0] n218_o;
  wire n220_o;
  wire [13:0] n221_o;
  reg [13:0] n222_o;
  wire [11:0] n223_o;
  wire [13:0] n225_o;
  wire [5:0] n226_o;
  wire [2:0] n227_o;
  wire [8:0] n228_o;
  wire [2:0] selfunctiontable4_n229;
  wire [2:0] selfunctiontable4_y;
  wire [13:0] n233_o;
  wire n235_o;
  wire n237_o;
  wire n238_o;
  wire [12:0] n240_o;
  wire [13:0] n242_o;
  wire n244_o;
  wire n246_o;
  wire n247_o;
  wire [1:0] n249_o;
  reg [13:0] n250_o;
  wire n251_o;
  wire [13:0] n252_o;
  wire n254_o;
  wire [13:0] n255_o;
  reg [13:0] n256_o;
  wire [11:0] n257_o;
  wire [13:0] n259_o;
  wire [5:0] n260_o;
  wire [2:0] n261_o;
  wire [8:0] n262_o;
  wire [2:0] selfunctiontable3_n263;
  wire [2:0] selfunctiontable3_y;
  wire [13:0] n267_o;
  wire n269_o;
  wire n271_o;
  wire n272_o;
  wire [12:0] n274_o;
  wire [13:0] n276_o;
  wire n278_o;
  wire n280_o;
  wire n281_o;
  wire [1:0] n283_o;
  reg [13:0] n284_o;
  wire n285_o;
  wire [13:0] n286_o;
  wire n288_o;
  wire [13:0] n289_o;
  reg [13:0] n290_o;
  wire [11:0] n291_o;
  wire [13:0] n293_o;
  wire [5:0] n294_o;
  wire [2:0] n295_o;
  wire [8:0] n296_o;
  wire [2:0] selfunctiontable2_n297;
  wire [2:0] selfunctiontable2_y;
  wire [13:0] n301_o;
  wire n303_o;
  wire n305_o;
  wire n306_o;
  wire [12:0] n308_o;
  wire [13:0] n310_o;
  wire n312_o;
  wire n314_o;
  wire n315_o;
  wire [1:0] n317_o;
  reg [13:0] n318_o;
  wire n319_o;
  wire [13:0] n320_o;
  wire n322_o;
  wire [13:0] n323_o;
  reg [13:0] n324_o;
  wire [11:0] n325_o;
  wire [13:0] n327_o;
  wire [5:0] n328_o;
  wire [2:0] n329_o;
  wire [8:0] n330_o;
  wire [2:0] selfunctiontable1_n331;
  wire [2:0] selfunctiontable1_y;
  wire [13:0] n335_o;
  wire n337_o;
  wire n339_o;
  wire n340_o;
  wire [12:0] n342_o;
  wire [13:0] n344_o;
  wire n346_o;
  wire n348_o;
  wire n349_o;
  wire [1:0] n351_o;
  reg [13:0] n352_o;
  wire n353_o;
  wire [13:0] n354_o;
  wire n356_o;
  wire [13:0] n357_o;
  reg [13:0] n358_o;
  wire [11:0] n359_o;
  wire n360_o;
  wire [1:0] n361_o;
  wire n362_o;
  wire [1:0] n364_o;
  wire [1:0] n365_o;
  wire n366_o;
  wire [1:0] n368_o;
  wire [1:0] n369_o;
  wire n370_o;
  wire [1:0] n372_o;
  wire [1:0] n373_o;
  wire n374_o;
  wire [1:0] n376_o;
  wire [1:0] n377_o;
  wire n378_o;
  wire [1:0] n380_o;
  wire [1:0] n381_o;
  wire n382_o;
  wire [1:0] n384_o;
  wire [1:0] n385_o;
  wire n386_o;
  wire [1:0] n388_o;
  wire [3:0] n389_o;
  wire [5:0] n390_o;
  wire [7:0] n391_o;
  wire [9:0] n392_o;
  wire [11:0] n393_o;
  wire [13:0] n394_o;
  wire n395_o;
  wire [2:0] n396_o;
  wire [4:0] n397_o;
  wire [6:0] n398_o;
  wire [8:0] n399_o;
  wire [10:0] n400_o;
  wire [12:0] n401_o;
  wire [13:0] n402_o;
  wire [13:0] n403_o;
  wire [12:0] n404_o;
  wire [10:0] n405_o;
  wire n406_o;
  wire [10:0] n407_o;
  wire [10:0] n408_o;
  wire n409_o;
  wire n410_o;
  wire [5:0] n412_o;
  wire [5:0] n413_o;
  wire [9:0] n414_o;
  wire [15:0] n415_o;
  wire [15:0] n417_o;
  wire [15:0] n418_o;
  wire n420_o;
  wire [1:0] n421_o;
  wire [1:0] n423_o;
  wire n425_o;
  wire [1:0] n426_o;
  wire n429_o;
  reg [1:0] n430_o;
  wire [2:0] n431_o;
  wire [13:0] n432_o;
  wire [16:0] n433_o;
  reg [5:0] n434_q;
  reg [5:0] n435_q;
  reg [5:0] n436_q;
  reg [5:0] n437_q;
  reg [5:0] n438_q;
  reg [5:0] n439_q;
  reg n440_q;
  reg n441_q;
  reg n442_q;
  reg n443_q;
  reg n444_q;
  reg n445_q;
  reg [1:0] n446_q;
  reg [1:0] n447_q;
  reg [1:0] n448_q;
  reg [1:0] n449_q;
  reg [1:0] n450_q;
  reg [1:0] n451_q;
  reg [10:0] n452_q;
  reg [10:0] n453_q;
  reg [10:0] n454_q;
  reg [10:0] n455_q;
  reg [10:0] n456_q;
  reg [13:0] n457_q;
  reg [2:0] n458_q;
  reg [13:0] n459_q;
  reg [2:0] n460_q;
  reg [13:0] n461_q;
  reg [2:0] n462_q;
  reg [13:0] n463_q;
  reg [13:0] n464_q;
  reg [2:0] n465_q;
  reg [13:0] n466_q;
  reg [13:0] n467_q;
  reg [2:0] n468_q;
  reg [1:0] n469_q;
  reg [1:0] n470_q;
  reg [1:0] n471_q;
  reg [1:0] n472_q;
  reg [1:0] n473_q;
  reg [1:0] n474_q;
  reg [1:0] n475_q;
  reg [1:0] n476_q;
  reg [1:0] n477_q;
  reg [1:0] n478_q;
  reg [1:0] n479_q;
  reg [1:0] n480_q;
  reg [1:0] n481_q;
  reg [1:0] n482_q;
  reg [1:0] n483_q;
  reg [1:0] n484_q;
  reg [1:0] n485_q;
  reg [1:0] n486_q;
  reg [1:0] n487_q;
  reg [1:0] n488_q;
  reg [1:0] n489_q;
  reg [1:0] n490_q;
  reg [1:0] n491_q;
  reg [1:0] n492_q;
  reg [1:0] n493_q;
  reg [1:0] n494_q;
  reg [1:0] n495_q;
  reg [1:0] n496_q;
  reg [1:0] n497_q;
  reg [1:0] n498_q;
  reg [1:0] n499_q;
  reg [1:0] n500_q;
  reg [1:0] n501_q;
  reg [1:0] n502_q;
  reg [1:0] n503_q;
  reg [1:0] n504_q;
  reg [13:0] n505_q;
  assign R = n433_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:588:8  */
  assign fx = n79_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:589:8  */
  assign fy = n82_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:8  */
  assign expr0 = n89_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:15  */
  assign expr0_d1 = n434_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:25  */
  assign expr0_d2 = n435_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:35  */
  assign expr0_d3 = n436_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:45  */
  assign expr0_d4 = n437_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:55  */
  assign expr0_d5 = n438_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:590:65  */
  assign expr0_d6 = n439_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:8  */
  assign sr = n92_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:12  */
  assign sr_d1 = n440_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:19  */
  assign sr_d2 = n441_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:26  */
  assign sr_d3 = n442_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:33  */
  assign sr_d4 = n443_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:40  */
  assign sr_d5 = n444_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:591:47  */
  assign sr_d6 = n445_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:592:8  */
  assign exnxy = n95_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:8  */
  assign exnr0 = n119_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:15  */
  assign exnr0_d1 = n446_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:25  */
  assign exnr0_d2 = n447_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:35  */
  assign exnr0_d3 = n448_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:45  */
  assign exnr0_d4 = n449_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:55  */
  assign exnr0_d5 = n450_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:593:65  */
  assign exnr0_d6 = n451_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:8  */
  assign d = fy; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:11  */
  assign d_d1 = n452_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:17  */
  assign d_d2 = n453_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:23  */
  assign d_d3 = n454_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:29  */
  assign d_d4 = n455_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:594:35  */
  assign d_d5 = n456_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:595:8  */
  assign psx = n121_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:596:8  */
  assign betaw7 = n123_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:597:8  */
  assign sel7 = n126_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:598:8  */
  assign q7 = q7_copy5; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:599:8  */
  assign q7_copy5 = selfunctiontable7_n127; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:600:8  */
  assign absq7d = n148_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:601:8  */
  assign w6 = n154_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:602:8  */
  assign betaw6 = n157_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:602:16  */
  assign betaw6_d1 = n457_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:603:8  */
  assign sel6 = n160_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:604:8  */
  assign q6 = q6_copy6_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:605:8  */
  assign q6_copy6 = selfunctiontable6_n161; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:605:18  */
  assign q6_copy6_d1 = n458_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:606:8  */
  assign absq6d = n182_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:607:8  */
  assign w5 = n188_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:608:8  */
  assign betaw5 = n191_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:608:16  */
  assign betaw5_d1 = n459_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:609:8  */
  assign sel5 = n194_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:610:8  */
  assign q5 = q5_copy7_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:611:8  */
  assign q5_copy7 = selfunctiontable5_n195; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:611:18  */
  assign q5_copy7_d1 = n460_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:612:8  */
  assign absq5d = n216_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:613:8  */
  assign w4 = n222_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:614:8  */
  assign betaw4 = n225_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:614:16  */
  assign betaw4_d1 = n461_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:615:8  */
  assign sel4 = n228_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:616:8  */
  assign q4 = q4_copy8; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:616:12  */
  assign q4_d1 = n462_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:617:8  */
  assign q4_copy8 = selfunctiontable4_n229; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:618:8  */
  assign absq4d = n250_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:618:16  */
  assign absq4d_d1 = n463_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:619:8  */
  assign w3 = n256_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:620:8  */
  assign betaw3 = n259_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:620:16  */
  assign betaw3_d1 = n464_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:621:8  */
  assign sel3 = n262_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:622:8  */
  assign q3 = q3_copy9; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:622:12  */
  assign q3_d1 = n465_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:623:8  */
  assign q3_copy9 = selfunctiontable3_n263; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:624:8  */
  assign absq3d = n284_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:624:16  */
  assign absq3d_d1 = n466_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:625:8  */
  assign w2 = n290_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:626:8  */
  assign betaw2 = n293_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:627:8  */
  assign sel2 = n296_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:628:8  */
  assign q2 = q2_copy10; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:629:8  */
  assign q2_copy10 = selfunctiontable2_n297; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:630:8  */
  assign absq2d = n318_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:631:8  */
  assign w1 = n324_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:632:8  */
  assign betaw1 = n327_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:632:16  */
  assign betaw1_d1 = n467_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:633:8  */
  assign sel1 = n330_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:634:8  */
  assign q1 = q1_copy11_d1; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:635:8  */
  assign q1_copy11 = selfunctiontable1_n331; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:635:19  */
  assign q1_copy11_d1 = n468_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:636:8  */
  assign absq1d = n352_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:637:8  */
  assign w0 = n358_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:638:8  */
  assign wfinal = n359_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:639:8  */
  assign qm0 = n360_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:8  */
  assign qp7 = n361_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:13  */
  assign qp7_d1 = n469_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:21  */
  assign qp7_d2 = n470_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:29  */
  assign qp7_d3 = n471_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:37  */
  assign qp7_d4 = n472_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:640:45  */
  assign qp7_d5 = n473_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:8  */
  assign qm7 = n364_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:13  */
  assign qm7_d1 = n474_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:21  */
  assign qm7_d2 = n475_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:29  */
  assign qm7_d3 = n476_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:37  */
  assign qm7_d4 = n477_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:641:45  */
  assign qm7_d5 = n478_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:642:8  */
  assign qp6 = n365_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:642:13  */
  assign qp6_d1 = n479_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:642:21  */
  assign qp6_d2 = n480_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:642:29  */
  assign qp6_d3 = n481_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:642:37  */
  assign qp6_d4 = n482_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:643:8  */
  assign qm6 = n368_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:643:13  */
  assign qm6_d1 = n483_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:643:21  */
  assign qm6_d2 = n484_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:643:29  */
  assign qm6_d3 = n485_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:643:37  */
  assign qm6_d4 = n486_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:644:8  */
  assign qp5 = n369_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:644:13  */
  assign qp5_d1 = n487_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:644:21  */
  assign qp5_d2 = n488_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:644:29  */
  assign qp5_d3 = n489_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:645:8  */
  assign qm5 = n372_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:645:13  */
  assign qm5_d1 = n490_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:645:21  */
  assign qm5_d2 = n491_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:645:29  */
  assign qm5_d3 = n492_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:646:8  */
  assign qp4 = n373_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:646:13  */
  assign qp4_d1 = n493_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:646:21  */
  assign qp4_d2 = n494_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:646:29  */
  assign qp4_d3 = n495_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:647:8  */
  assign qm4 = n376_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:647:13  */
  assign qm4_d1 = n496_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:647:21  */
  assign qm4_d2 = n497_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:647:29  */
  assign qm4_d3 = n498_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:648:8  */
  assign qp3 = n377_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:648:13  */
  assign qp3_d1 = n499_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:648:21  */
  assign qp3_d2 = n500_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:649:8  */
  assign qm3 = n380_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:649:13  */
  assign qm3_d1 = n501_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:649:21  */
  assign qm3_d2 = n502_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:650:8  */
  assign qp2 = n381_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:650:13  */
  assign qp2_d1 = n503_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:651:8  */
  assign qm2 = n384_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:651:13  */
  assign qm2_d1 = n504_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:652:8  */
  assign qp1 = n385_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:653:8  */
  assign qm1 = n388_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:654:8  */
  assign qp = n394_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:655:8  */
  assign qm = n402_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:656:8  */
  assign quotient = n403_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:656:18  */
  assign quotient_d1 = n505_q; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:657:8  */
  assign mr = n404_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:658:8  */
  assign frnorm = n407_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:659:8  */
  assign round = n409_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:660:8  */
  assign expr1 = n413_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:661:8  */
  assign expfrac = n415_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:662:8  */
  assign expfracr = n418_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:663:8  */
  assign exnr = n421_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:664:8  */
  assign exnrfinal = n430_o; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:743:17  */
  assign n77_o = X[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:743:14  */
  assign n79_o = {1'b1, n77_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:744:17  */
  assign n80_o = Y[9:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:744:14  */
  assign n82_o = {1'b1, n80_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:746:22  */
  assign n83_o = X[13:10];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:746:19  */
  assign n85_o = {2'b00, n83_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:746:49  */
  assign n86_o = Y[13:10];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:746:46  */
  assign n88_o = {2'b00, n86_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:746:38  */
  assign n89_o = n85_o - n88_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:747:11  */
  assign n90_o = X[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:747:21  */
  assign n91_o = Y[14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:747:16  */
  assign n92_o = n90_o ^ n91_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:749:14  */
  assign n93_o = X[16:15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:749:32  */
  assign n94_o = Y[16:15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:749:29  */
  assign n95_o = {n93_o, n94_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:752:18  */
  assign n98_o = exnxy == 4'b0101;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:753:18  */
  assign n101_o = exnxy == 4'b0001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:753:30  */
  assign n103_o = exnxy == 4'b0010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:753:30  */
  assign n104_o = n101_o | n103_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:753:39  */
  assign n106_o = exnxy == 4'b0110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:753:39  */
  assign n107_o = n104_o | n106_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:754:18  */
  assign n110_o = exnxy == 4'b0100;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:754:30  */
  assign n112_o = exnxy == 4'b1000;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:754:30  */
  assign n113_o = n110_o | n112_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:754:39  */
  assign n115_o = exnxy == 4'b1001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:754:39  */
  assign n116_o = n113_o | n115_o;
  assign n118_o = {n116_o, n107_o, n98_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:750:4  */
  always @*
    case (n118_o)
      3'b100: n119_o = 2'b10;
      3'b010: n119_o = 2'b00;
      3'b001: n119_o = 2'b01;
      default: n119_o = 2'b11;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:757:15  */
  assign n121_o = {1'b0, fx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:758:20  */
  assign n123_o = {2'b00, psx};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:759:18  */
  assign n124_o = betaw7[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:759:35  */
  assign n125_o = d[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:759:32  */
  assign n126_o = {n124_o, n125_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:762:23  */
  assign selfunctiontable7_n127 = selfunctiontable7_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:760:4  */
  selfunction_f300_uid4 selfunctiontable7 (
    .x(sel7),
    .y(selfunctiontable7_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:767:16  */
  assign n131_o = {3'b000, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:767:66  */
  assign n133_o = q7 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:767:77  */
  assign n135_o = q7 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:767:77  */
  assign n136_o = n133_o | n135_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:768:15  */
  assign n138_o = {2'b00, d};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:768:19  */
  assign n140_o = {n138_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:768:52  */
  assign n142_o = q7 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:768:63  */
  assign n144_o = q7 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:768:63  */
  assign n145_o = n142_o | n144_o;
  assign n147_o = {n145_o, n136_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:765:4  */
  always @*
    case (n147_o)
      2'b10: n148_o = n140_o;
      2'b01: n148_o = n131_o;
      default: n148_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:771:11  */
  assign n149_o = q7[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:772:16  */
  assign n150_o = betaw7 - absq7d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:772:25  */
  assign n152_o = n149_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:773:17  */
  assign n153_o = betaw7 + absq7d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:771:4  */
  always @*
    case (n152_o)
      1'b1: n154_o = n150_o;
      default: n154_o = n153_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:775:16  */
  assign n155_o = w6[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:775:30  */
  assign n157_o = {n155_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:776:18  */
  assign n158_o = betaw6[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:776:35  */
  assign n159_o = d[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:776:32  */
  assign n160_o = {n158_o, n159_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:779:23  */
  assign selfunctiontable6_n161 = selfunctiontable6_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:777:4  */
  selfunction_f300_uid4 selfunctiontable6 (
    .x(sel6),
    .y(selfunctiontable6_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:784:16  */
  assign n165_o = {3'b000, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:784:66  */
  assign n167_o = q6 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:784:77  */
  assign n169_o = q6 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:784:77  */
  assign n170_o = n167_o | n169_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:785:15  */
  assign n172_o = {2'b00, d_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:785:22  */
  assign n174_o = {n172_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:785:52  */
  assign n176_o = q6 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:785:63  */
  assign n178_o = q6 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:785:63  */
  assign n179_o = n176_o | n178_o;
  assign n181_o = {n179_o, n170_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:782:4  */
  always @*
    case (n181_o)
      2'b10: n182_o = n174_o;
      2'b01: n182_o = n165_o;
      default: n182_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:788:11  */
  assign n183_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:789:19  */
  assign n184_o = betaw6_d1 - absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:789:28  */
  assign n186_o = n183_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:790:20  */
  assign n187_o = betaw6_d1 + absq6d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:788:4  */
  always @*
    case (n186_o)
      1'b1: n188_o = n184_o;
      default: n188_o = n187_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:792:16  */
  assign n189_o = w5[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:792:30  */
  assign n191_o = {n189_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:793:18  */
  assign n192_o = betaw5[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:793:38  */
  assign n193_o = d_d1[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:793:32  */
  assign n194_o = {n192_o, n193_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:796:23  */
  assign selfunctiontable5_n195 = selfunctiontable5_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:794:4  */
  selfunction_f300_uid4 selfunctiontable5 (
    .x(sel5),
    .y(selfunctiontable5_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:801:16  */
  assign n199_o = {3'b000, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:801:66  */
  assign n201_o = q5 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:801:77  */
  assign n203_o = q5 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:801:77  */
  assign n204_o = n201_o | n203_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:802:15  */
  assign n206_o = {2'b00, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:802:22  */
  assign n208_o = {n206_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:802:52  */
  assign n210_o = q5 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:802:63  */
  assign n212_o = q5 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:802:63  */
  assign n213_o = n210_o | n212_o;
  assign n215_o = {n213_o, n204_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:799:4  */
  always @*
    case (n215_o)
      2'b10: n216_o = n208_o;
      2'b01: n216_o = n199_o;
      default: n216_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:805:11  */
  assign n217_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:806:19  */
  assign n218_o = betaw5_d1 - absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:806:28  */
  assign n220_o = n217_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:807:20  */
  assign n221_o = betaw5_d1 + absq5d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:805:4  */
  always @*
    case (n220_o)
      1'b1: n222_o = n218_o;
      default: n222_o = n221_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:809:16  */
  assign n223_o = w4[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:809:30  */
  assign n225_o = {n223_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:810:18  */
  assign n226_o = betaw4[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:810:38  */
  assign n227_o = d_d2[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:810:32  */
  assign n228_o = {n226_o, n227_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:813:23  */
  assign selfunctiontable4_n229 = selfunctiontable4_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:811:4  */
  selfunction_f300_uid4 selfunctiontable4 (
    .x(sel4),
    .y(selfunctiontable4_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:818:16  */
  assign n233_o = {3'b000, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:818:66  */
  assign n235_o = q4 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:818:77  */
  assign n237_o = q4 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:818:77  */
  assign n238_o = n235_o | n237_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:819:15  */
  assign n240_o = {2'b00, d_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:819:22  */
  assign n242_o = {n240_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:819:52  */
  assign n244_o = q4 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:819:63  */
  assign n246_o = q4 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:819:63  */
  assign n247_o = n244_o | n246_o;
  assign n249_o = {n247_o, n238_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:816:4  */
  always @*
    case (n249_o)
      2'b10: n250_o = n242_o;
      2'b01: n250_o = n233_o;
      default: n250_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:822:14  */
  assign n251_o = q4_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:823:19  */
  assign n252_o = betaw4_d1 - absq4d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:823:31  */
  assign n254_o = n251_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:824:20  */
  assign n255_o = betaw4_d1 + absq4d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:822:4  */
  always @*
    case (n254_o)
      1'b1: n256_o = n252_o;
      default: n256_o = n255_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:826:16  */
  assign n257_o = w3[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:826:30  */
  assign n259_o = {n257_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:827:18  */
  assign n260_o = betaw3[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:827:38  */
  assign n261_o = d_d3[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:827:32  */
  assign n262_o = {n260_o, n261_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:830:23  */
  assign selfunctiontable3_n263 = selfunctiontable3_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:828:4  */
  selfunction_f300_uid4 selfunctiontable3 (
    .x(sel3),
    .y(selfunctiontable3_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:835:16  */
  assign n267_o = {3'b000, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:835:66  */
  assign n269_o = q3 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:835:77  */
  assign n271_o = q3 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:835:77  */
  assign n272_o = n269_o | n271_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:836:15  */
  assign n274_o = {2'b00, d_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:836:22  */
  assign n276_o = {n274_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:836:52  */
  assign n278_o = q3 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:836:63  */
  assign n280_o = q3 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:836:63  */
  assign n281_o = n278_o | n280_o;
  assign n283_o = {n281_o, n272_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:833:4  */
  always @*
    case (n283_o)
      2'b10: n284_o = n276_o;
      2'b01: n284_o = n267_o;
      default: n284_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:839:14  */
  assign n285_o = q3_d1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:840:19  */
  assign n286_o = betaw3_d1 - absq3d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:840:31  */
  assign n288_o = n285_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:841:20  */
  assign n289_o = betaw3_d1 + absq3d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:839:4  */
  always @*
    case (n288_o)
      1'b1: n290_o = n286_o;
      default: n290_o = n289_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:843:16  */
  assign n291_o = w2[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:843:30  */
  assign n293_o = {n291_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:844:18  */
  assign n294_o = betaw2[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:844:38  */
  assign n295_o = d_d4[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:844:32  */
  assign n296_o = {n294_o, n295_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:847:23  */
  assign selfunctiontable2_n297 = selfunctiontable2_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:845:4  */
  selfunction_f300_uid4 selfunctiontable2 (
    .x(sel2),
    .y(selfunctiontable2_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:852:16  */
  assign n301_o = {3'b000, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:852:66  */
  assign n303_o = q2 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:852:77  */
  assign n305_o = q2 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:852:77  */
  assign n306_o = n303_o | n305_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:853:15  */
  assign n308_o = {2'b00, d_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:853:22  */
  assign n310_o = {n308_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:853:52  */
  assign n312_o = q2 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:853:63  */
  assign n314_o = q2 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:853:63  */
  assign n315_o = n312_o | n314_o;
  assign n317_o = {n315_o, n306_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:850:4  */
  always @*
    case (n317_o)
      2'b10: n318_o = n310_o;
      2'b01: n318_o = n301_o;
      default: n318_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:856:11  */
  assign n319_o = q2[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:857:16  */
  assign n320_o = betaw2 - absq2d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:857:25  */
  assign n322_o = n319_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:858:17  */
  assign n323_o = betaw2 + absq2d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:856:4  */
  always @*
    case (n322_o)
      1'b1: n324_o = n320_o;
      default: n324_o = n323_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:860:16  */
  assign n325_o = w1[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:860:30  */
  assign n327_o = {n325_o, 2'b00};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:861:18  */
  assign n328_o = betaw1[13:8];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:861:38  */
  assign n329_o = d_d4[9:7];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:861:32  */
  assign n330_o = {n328_o, n329_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:864:23  */
  assign selfunctiontable1_n331 = selfunctiontable1_y; // (signal)
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:862:4  */
  selfunction_f300_uid4 selfunctiontable1 (
    .x(sel1),
    .y(selfunctiontable1_y));
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:869:16  */
  assign n335_o = {3'b000, d_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:869:66  */
  assign n337_o = q1 == 3'b001;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:869:77  */
  assign n339_o = q1 == 3'b111;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:869:77  */
  assign n340_o = n337_o | n339_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:870:15  */
  assign n342_o = {2'b00, d_d5};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:870:22  */
  assign n344_o = {n342_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:870:52  */
  assign n346_o = q1 == 3'b010;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:870:63  */
  assign n348_o = q1 == 3'b110;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:870:63  */
  assign n349_o = n346_o | n348_o;
  assign n351_o = {n349_o, n340_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:867:4  */
  always @*
    case (n351_o)
      2'b10: n352_o = n344_o;
      2'b01: n352_o = n335_o;
      default: n352_o = 14'b00000000000000;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:873:11  */
  assign n353_o = q1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:874:19  */
  assign n354_o = betaw1_d1 - absq1d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:874:28  */
  assign n356_o = n353_o == 1'b0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:875:20  */
  assign n357_o = betaw1_d1 + absq1d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:873:4  */
  always @*
    case (n356_o)
      1'b1: n358_o = n354_o;
      default: n358_o = n357_o;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:877:16  */
  assign n359_o = w0[11:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:878:17  */
  assign n360_o = wfinal[11];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:879:18  */
  assign n361_o = q7[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:880:18  */
  assign n362_o = q7[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:880:22  */
  assign n364_o = {n362_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:881:18  */
  assign n365_o = q6[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:882:18  */
  assign n366_o = q6[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:882:22  */
  assign n368_o = {n366_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:883:18  */
  assign n369_o = q5[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:884:18  */
  assign n370_o = q5[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:884:22  */
  assign n372_o = {n370_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:885:18  */
  assign n373_o = q4[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:886:18  */
  assign n374_o = q4[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:886:22  */
  assign n376_o = {n374_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:887:18  */
  assign n377_o = q3[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:888:18  */
  assign n378_o = q3[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:888:22  */
  assign n380_o = {n378_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:889:18  */
  assign n381_o = q2[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:890:18  */
  assign n382_o = q2[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:890:22  */
  assign n384_o = {n382_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:891:18  */
  assign n385_o = q1[1:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:892:18  */
  assign n386_o = q1[2];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:892:22  */
  assign n388_o = {n386_o, 1'b0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:17  */
  assign n389_o = {qp7_d5, qp6_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:26  */
  assign n390_o = {n389_o, qp5_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:35  */
  assign n391_o = {n390_o, qp4_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:44  */
  assign n392_o = {n391_o, qp3_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:53  */
  assign n393_o = {n392_o, qp2_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:893:62  */
  assign n394_o = {n393_o, qp1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:16  */
  assign n395_o = qm7_d5[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:20  */
  assign n396_o = {n395_o, qm6_d4};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:29  */
  assign n397_o = {n396_o, qm5_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:38  */
  assign n398_o = {n397_o, qm4_d3};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:47  */
  assign n399_o = {n398_o, qm3_d2};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:56  */
  assign n400_o = {n399_o, qm2_d1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:65  */
  assign n401_o = {n400_o, qm1};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:894:71  */
  assign n402_o = {n401_o, qm0};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:895:19  */
  assign n403_o = qp - qm;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:899:21  */
  assign n404_o = quotient_d1[12:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:901:19  */
  assign n405_o = mr[11:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:901:41  */
  assign n406_o = mr[12];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:901:34  */
  assign n407_o = n406_o ? n405_o : n408_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:902:19  */
  assign n408_o = mr[10:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:903:19  */
  assign n409_o = frnorm[0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:904:57  */
  assign n410_o = mr[12];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:904:53  */
  assign n412_o = {5'b00011, n410_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:904:22  */
  assign n413_o = expr0_d6 + n412_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:906:29  */
  assign n414_o = frnorm[10:1];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:906:21  */
  assign n415_o = {expr1, n414_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:907:48  */
  assign n417_o = {15'b000000000000000, round};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:907:24  */
  assign n418_o = expfrac + n417_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:908:36  */
  assign n420_o = expfracr[15];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:908:23  */
  assign n421_o = n420_o ? 2'b00 : n426_o;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:909:37  */
  assign n423_o = expfracr[15:14];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:909:52  */
  assign n425_o = n423_o == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:909:12  */
  assign n426_o = n425_o ? 2'b10 : 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:913:17  */
  assign n429_o = exnr0_d6 == 2'b01;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:911:4  */
  always @*
    case (n429_o)
      1'b1: n430_o = exnr;
      default: n430_o = exnr0_d6;
    endcase
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:915:19  */
  assign n431_o = {exnrfinal, sr_d6};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:915:37  */
  assign n432_o = expfracr[13:0];
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:915:27  */
  assign n433_o = {n431_o, n432_o};
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n434_q <= expr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n435_q <= expr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n436_q <= expr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n437_q <= expr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n438_q <= expr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n439_q <= expr0_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n440_q <= sr;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n441_q <= sr_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n442_q <= sr_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n443_q <= sr_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n444_q <= sr_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n445_q <= sr_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n446_q <= exnr0;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n447_q <= exnr0_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n448_q <= exnr0_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n449_q <= exnr0_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n450_q <= exnr0_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n451_q <= exnr0_d5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n452_q <= d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n453_q <= d_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n454_q <= d_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n455_q <= d_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n456_q <= d_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n457_q <= betaw6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n458_q <= q6_copy6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n459_q <= betaw5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n460_q <= q5_copy7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n461_q <= betaw4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n462_q <= q4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n463_q <= absq4d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n464_q <= betaw3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n465_q <= q3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n466_q <= absq3d;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n467_q <= betaw1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n468_q <= q1_copy11;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n469_q <= qp7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n470_q <= qp7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n471_q <= qp7_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n472_q <= qp7_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n473_q <= qp7_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n474_q <= qm7;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n475_q <= qm7_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n476_q <= qm7_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n477_q <= qm7_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n478_q <= qm7_d4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n479_q <= qp6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n480_q <= qp6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n481_q <= qp6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n482_q <= qp6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n483_q <= qm6;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n484_q <= qm6_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n485_q <= qm6_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n486_q <= qm6_d3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n487_q <= qp5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n488_q <= qp5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n489_q <= qp5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n490_q <= qm5;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n491_q <= qm5_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n492_q <= qm5_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n493_q <= qp4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n494_q <= qp4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n495_q <= qp4_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n496_q <= qm4;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n497_q <= qm4_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n498_q <= qm4_d2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n499_q <= qp3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n500_q <= qp3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n501_q <= qm3;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n502_q <= qm3_d1;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n503_q <= qp2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n504_q <= qm2;
  /* /home/mlevental/dev_projects/bragghls/scripts/../bragghls/ip_cores/flopoco_fdiv_4_10.vhdl:668:10  */
  always @(posedge clk)
    n505_q <= quotient;
endmodule

